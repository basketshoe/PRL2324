library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity Test_8214 is
end Test_8214;

architecture ARCH of Test_8214 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

	signal memory_control : std_logic := '0';
	
	signal continue : std_logic := '0';

-- Scenario Definition

	--Scenario 0
	constant SCENARIO_LENGTH_0 : integer := 1020;
	type scenario_type_0 is array (0 to SCENARIO_LENGTH_0*2-1) of integer;
	signal scenario_input_0 : scenario_type_0 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 100,   0, 137,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 151,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  85,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 209,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 111,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 111,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 163,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  48,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 191,   0,   0,   0, 122,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  23,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 212,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  20,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 176,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 189,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 224,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 190,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 209,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 175,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  88,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 106,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 119,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 242,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  67,   0,   0,   0,   0,   0,   0,   0, 113,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  63,   0,   0,   0,   0,   0,   0,   0,  50,   0,   0,   0,   0,   0,   0,   0,   0,   0, 118,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_0  : scenario_type_0 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 100,  31, 137,  31, 137,  30, 137,  29, 137,  28, 137,  27, 137,  26, 137,  25, 137,  24, 137,  23, 137,  22, 137,  21, 137,  20, 137,  19, 137,  18, 137,  17, 137,  16, 137,  15, 137,  14, 137,  13, 137,  12, 137,  11, 137,  10, 137,   9, 137,   8, 137,   7, 137,   6, 137,   5, 137,   4, 137,   3, 137,   2, 137,   1, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 151,  31, 151,  30, 151,  29, 151,  28, 151,  27, 151,  26, 151,  25, 151,  24, 151,  23, 151,  22, 151,  21, 151,  20, 151,  19, 151,  18, 151,  17, 151,  16, 151,  15, 151,  14, 151,  13, 151,  12, 151,  11, 151,  10, 151,   9, 151,   8, 151,   7, 151,   6, 151,   5, 151,   4, 151,   3, 151,   2, 151,   1, 151,   0, 151,   0, 151,   0, 151,   0, 151,   0, 151,   0, 151,   0, 151,   0, 151,   0, 151,   0, 151,   0, 151,   0, 151,   0,  85,  31,  85,  30,  85,  29,  85,  28,  85,  27,  85,  26,  85,  25,  85,  24,  85,  23,  85,  22,  85,  21,  85,  20,  85,  19,  85,  18,  85,  17,  85,  16,  85,  15,  85,  14,  85,  13,  85,  12,  85,  11,  85,  10,  85,   9,  85,   8,  85,   7,  85,   6,  85,   5,  85,   4,  85,   3,  85,   2, 209,  31, 209,  30, 209,  29, 209,  28, 209,  27, 209,  26, 209,  25, 209,  24, 209,  23, 209,  22, 209,  21, 209,  20, 209,  19, 209,  18, 209,  17, 209,  16, 209,  15, 209,  14, 209,  13, 111,  31, 111,  30, 111,  29, 111,  28, 111,  27, 111,  26, 111,  25, 111,  24, 111,  23, 111,  22, 111,  21, 111,  31, 111,  30, 111,  29, 111,  28, 111,  27, 111,  26, 111,  25, 111,  24, 111,  23, 111,  22, 111,  21, 111,  20, 111,  19, 111,  18, 111,  17, 111,  16, 111,  15, 111,  14, 111,  13, 111,  12, 111,  11, 111,  10, 111,   9, 111,   8, 111,   7, 111,   6, 111,   5, 111,   4, 111,   3, 111,   2, 111,   1, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 163,  31, 163,  30, 163,  29, 163,  28, 163,  27, 163,  26, 163,  25, 163,  24, 163,  23, 163,  22, 163,  21, 163,  20, 163,  19, 163,  18, 163,  17, 163,  16, 163,  15, 163,  14, 163,  13, 163,  12, 163,  11, 163,  10, 163,   9, 163,   8,  48,  31,  48,  30,  48,  29,  48,  28,  48,  27,  48,  26,  48,  25,  48,  24,  48,  23,  48,  22,  48,  21,  48,  20,  48,  19,  48,  18,  48,  17,  48,  16,  48,  15,  48,  14,  48,  13,  48,  12,  48,  11,  48,  10,  48,   9,  48,   8,  48,   7,  48,   6,  48,   5,  48,   4,  48,   3,  48,   2,  48,   1,  48,   0,  48,   0,  48,   0,  48,   0,  48,   0,  48,   0,  48,   0,  48,   0,  48,   0,  48,   0,  48,   0,  48,   0,  48,   0,  48,   0,  48,   0,  48,   0,  48,   0, 191,  31, 191,  30, 122,  31, 122,  30, 122,  29, 122,  28, 122,  27, 122,  26, 122,  25, 122,  24, 122,  23, 122,  22, 122,  21, 122,  20, 122,  19, 122,  18, 122,  17, 122,  16, 122,  15, 122,  14, 122,  13, 122,  12, 122,  11, 122,  10, 122,   9,  23,  31,  23,  30,  23,  29,  23,  28,  23,  27,  23,  26,  23,  25,  23,  24,  23,  23,  23,  22,  23,  21,  23,  20,  23,  19,  23,  18,  23,  17,  23,  16,  23,  15,  23,  14,  23,  13,  23,  12,  23,  11,  23,  10,  23,   9,  23,   8,  23,   7,  23,   6,  23,   5,  23,   4,  23,   3,  23,   2,  23,   1,  23,   0,  23,   0,  23,   0,  23,   0,  23,   0,  23,   0,  23,   0,  23,   0,  23,   0,  23,   0,  23,   0,  23,   0, 212,  31, 212,  30, 212,  29, 212,  28, 212,  27, 212,  26, 212,  25, 212,  24, 212,  23, 212,  22, 212,  21, 212,  20, 212,  19, 212,  18, 212,  17, 212,  16, 212,  15, 212,  14, 212,  13, 212,  12, 212,  11, 212,  10, 212,   9, 212,   8, 212,   7, 212,   6, 212,   5, 212,   4, 212,   3, 212,   2, 212,   1, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0,  20,  31,  20,  30,  20,  29,  20,  28,  20,  27,  20,  26,  20,  25,  20,  24,  20,  23,  20,  22,  20,  21,  20,  20,  20,  19,  20,  18,  20,  17,  20,  16,  20,  15,  20,  14,  20,  13,  20,  12,  20,  11,  20,  10,  20,   9,  20,   8, 176,  31, 176,  30, 176,  29, 176,  28, 176,  27, 176,  26, 176,  25, 176,  24, 176,  23, 176,  22, 176,  21, 176,  20, 176,  19, 176,  18, 176,  17, 176,  16, 176,  15, 176,  14, 176,  13, 176,  12, 189,  31, 189,  30, 189,  29, 189,  28, 189,  27, 189,  26, 189,  25, 189,  24, 189,  23, 189,  22, 189,  21, 189,  20, 189,  19, 189,  18, 189,  17, 189,  16, 189,  15, 189,  14, 189,  13, 189,  12, 189,  11, 189,  10, 189,   9, 189,   8, 189,   7, 189,   6, 189,   5, 189,   4, 189,   3, 189,   2, 189,   1, 189,   0, 189,   0, 189,   0, 189,   0, 189,   0, 224,  31, 224,  30, 224,  29, 224,  28, 224,  27, 224,  26, 224,  25, 224,  24, 224,  23, 190,  31, 190,  30, 190,  29, 190,  28, 190,  27, 190,  26, 190,  25, 190,  24, 190,  23, 190,  22, 190,  21, 190,  20, 190,  19, 190,  18, 209,  31, 209,  30, 209,  29, 209,  28, 209,  27, 209,  26, 209,  25, 209,  24, 209,  23, 209,  22, 209,  21, 209,  20, 209,  19, 209,  18, 209,  17, 209,  16, 209,  15, 209,  14, 209,  13, 209,  12, 209,  11, 209,  10, 175,  31, 175,  30, 175,  29, 175,  28, 175,  27, 175,  26, 175,  25, 175,  24, 175,  23, 175,  22, 175,  21, 175,  20, 175,  19, 175,  18, 175,  17, 175,  16, 175,  15, 175,  14, 175,  13, 175,  12, 175,  11, 175,  10, 175,   9, 175,   8, 175,   7, 175,   6, 175,   5, 175,   4, 175,   3, 175,   2, 175,   1, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0, 175,   0,  88,  31,  88,  30,  88,  29,  88,  28,  88,  27,  88,  26,  88,  25,  88,  24,  88,  23,  88,  22,  88,  21,  88,  20,  88,  19,  88,  18,  88,  17,  88,  16,  88,  15,  88,  14,  88,  13,  88,  12, 106,  31, 106,  30, 106,  29, 106,  28, 106,  27, 106,  26, 106,  25, 106,  24, 106,  23, 106,  22, 106,  21, 106,  20, 106,  19, 106,  18, 106,  17, 106,  16, 106,  15, 106,  14, 106,  13, 106,  12, 106,  11, 106,  10, 106,   9, 106,   8, 106,   7, 106,   6, 106,   5, 106,   4, 106,   3, 119,  31, 119,  30, 119,  29, 119,  28, 119,  27, 119,  26, 119,  25, 119,  24, 119,  23, 119,  22, 119,  21, 119,  20, 119,  19, 119,  18, 119,  17, 119,  16, 119,  15, 119,  14, 119,  13, 119,  12, 119,  11, 119,  10, 119,   9, 119,   8, 119,   7, 119,   6, 119,   5, 119,   4, 119,   3, 119,   2, 119,   1, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 242,  31, 242,  30, 242,  29, 242,  28, 242,  27, 242,  26, 242,  25, 242,  24, 242,  23, 242,  22, 242,  21, 242,  20,  67,  31,  67,  30,  67,  29,  67,  28, 113,  31, 113,  30, 113,  29, 113,  28, 113,  27, 113,  26, 113,  25, 113,  24, 113,  23, 113,  22, 113,  21, 113,  20, 113,  19, 113,  18, 113,  17, 113,  16, 113,  15, 113,  14, 113,  13, 113,  12, 113,  11, 113,  10, 113,   9, 113,   8, 113,   7, 113,   6, 113,   5, 113,   4, 113,   3, 113,   2, 113,   1, 113,   0, 113,   0, 113,   0, 113,   0, 113,   0, 113,   0, 113,   0,  63,  31,  63,  30,  63,  29,  63,  28,  50,  31,  50,  30,  50,  29,  50,  28,  50,  27, 118,  31, 118,  30, 118,  29, 118,  28, 118,  27, 118,  26, 118,  25, 118,  24, 118,  23, 118,  22, 118,  21, 118,  20, 118,  19, 118,  18, 118,  17, 118,  16, 118,  15, 118,  14, 118,  13, 118,  12, 118,  11, 118,  10, 118,   9, 118,   8, 118,   7, 118,   6, 118,   5);
	constant SCENARIO_ADDRESS_0 : integer := 7;


	--Scenario 1
	constant SCENARIO_LENGTH_1 : integer := 1019;
	type scenario_type_1 is array (0 to SCENARIO_LENGTH_1*2-1) of integer;
	signal scenario_input_1 : scenario_type_1 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 182,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  11,   0,   0,   0, 240,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 164,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  91,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 212,   0,   0,   0,   0,   0,   0,   0, 136,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 161,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 135,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  82,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  51,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  81,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 160,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 137,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   5,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 145,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  41,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 244,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 218,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 144,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  13,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 160,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 125,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_1  : scenario_type_1 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 182,  31, 182,  30, 182,  29, 182,  28, 182,  27, 182,  26, 182,  25, 182,  24, 182,  23, 182,  22, 182,  21, 182,  20, 182,  19, 182,  18, 182,  17, 182,  16, 182,  15, 182,  14, 182,  13, 182,  12, 182,  11, 182,  10, 182,   9, 182,   8, 182,   7, 182,   6, 182,   5, 182,   4, 182,   3, 182,   2, 182,   1, 182,   0, 182,   0, 182,   0, 182,   0, 182,   0, 182,   0, 182,   0, 182,   0, 182,   0, 182,   0,  11,  31,  11,  30, 240,  31, 240,  30, 240,  29, 240,  28, 240,  27, 240,  26, 240,  25, 240,  24, 240,  23, 240,  22, 240,  21, 240,  20, 240,  19, 240,  18, 240,  17, 240,  16, 240,  15, 240,  14, 240,  13, 240,  12, 240,  11, 240,  10, 240,   9, 240,   8, 240,   7, 240,   6, 240,   5, 240,   4, 240,   3, 240,   2, 240,   1, 240,   0, 240,   0, 240,   0, 240,   0, 240,   0, 240,   0, 240,   0, 240,   0, 240,   0, 240,   0, 240,   0, 240,   0, 240,   0, 240,   0, 240,   0, 240,   0, 164,  31, 164,  30, 164,  29, 164,  28, 164,  27, 164,  26, 164,  25, 164,  24, 164,  23, 164,  22, 164,  21, 164,  20, 164,  19, 164,  18, 164,  17, 164,  16, 164,  15, 164,  14, 164,  13, 164,  12, 164,  11, 164,  10, 164,   9, 164,   8, 164,   7, 164,   6, 164,   5, 164,   4, 164,   3, 164,   2,  91,  31,  91,  30,  91,  29,  91,  28,  91,  27,  91,  26,  91,  25,  91,  24,  91,  23,  91,  22,  91,  21,  91,  20,  91,  19,  91,  18,  91,  17,  91,  16,  91,  15,  91,  14,  91,  13,  91,  12,  91,  11,  91,  10,  91,   9,  91,   8,  91,   7,  91,   6,  91,   5,  91,   4,  91,   3,  91,   2,  91,   1,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0, 212,  31, 212,  30, 212,  29, 212,  28, 136,  31, 136,  30, 136,  29, 136,  28, 136,  27, 136,  26, 136,  25, 136,  24, 161,  31, 161,  30, 161,  29, 161,  28, 161,  27, 161,  26, 161,  25, 161,  24, 161,  23, 161,  22, 161,  21, 161,  20, 161,  19, 161,  18, 161,  17, 161,  16, 161,  15, 161,  14, 161,  13, 161,  12, 161,  11, 161,  10, 161,   9, 161,   8, 161,   7, 161,   6, 161,   5, 161,   4, 161,   3, 161,   2, 161,   1, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 135,  31, 135,  30, 135,  29, 135,  28, 135,  27, 135,  26, 135,  25, 135,  24, 135,  23, 135,  22, 135,  21, 135,  20, 135,  19, 135,  18, 135,  17,  82,  31,  82,  30,  82,  29,  82,  28,  82,  27,  82,  26,  82,  25,  82,  24,  82,  23,  82,  22,  82,  21,  82,  20,  82,  19,  82,  18,  82,  17,  82,  16,  82,  15,  82,  14,  82,  13,  82,  12,  82,  11,  82,  10,  82,   9,  82,   8,  82,   7,  82,   6,  82,   5,  82,   4,  82,   3,  82,   2,  82,   1,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  51,  31,  51,  30,  51,  29,  51,  28,  51,  27,  51,  26,  51,  25,  51,  24,  51,  23,  51,  22,  51,  21,  51,  20,  51,  19,  51,  18,  51,  17,  51,  16,  51,  15,  51,  14,  51,  13,  51,  12,  51,  11,  51,  10,  51,   9,  51,   8,  51,   7,  51,   6,  51,   5,  51,   4,  51,   3,  51,   2,  51,   1,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  81,  31,  81,  30,  81,  29,  81,  28,  81,  27,  81,  26,  81,  25,  81,  24,  81,  23,  81,  22,  81,  21,  81,  20,  81,  19,  81,  18,  81,  17,  81,  16,  81,  15,  81,  14,  81,  13,  81,  12,  81,  11,  81,  10,  81,   9,  81,   8,  81,   7,  81,   6,  81,   5,  81,   4,  81,   3,  81,   2,  81,   1,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0,  81,   0, 160,  31, 160,  30, 160,  29, 160,  28, 160,  27, 160,  26, 160,  25, 160,  24, 160,  23, 160,  22, 160,  21, 160,  20, 160,  19, 160,  18, 160,  17, 160,  16, 160,  15, 160,  14, 160,  13, 160,  12, 160,  11, 160,  10, 160,   9, 160,   8, 160,   7, 160,   6, 160,   5, 160,   4, 160,   3, 160,   2, 160,   1, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 137,  31, 137,  30, 137,  29, 137,  28, 137,  27, 137,  26, 137,  25, 137,  24, 137,  23, 137,  22, 137,  21, 137,  20, 137,  19, 137,  18, 137,  17, 137,  16, 137,  15, 137,  14, 137,  13, 137,  12, 137,  11, 137,  10, 137,   9, 137,   8, 137,   7, 137,   6,   5,  31,   5,  30,   5,  29,   5,  28,   5,  27,   5,  26,   5,  25,   5,  24,   5,  23,   5,  22,   5,  21,   5,  20, 145,  31, 145,  30, 145,  29, 145,  28, 145,  27, 145,  26, 145,  25, 145,  24, 145,  23, 145,  22, 145,  21, 145,  20, 145,  19, 145,  18, 145,  17, 145,  16, 145,  15, 145,  14, 145,  13, 145,  12, 145,  11, 145,  10, 145,   9, 145,   8, 145,   7, 145,   6, 145,   5, 145,   4, 145,   3, 145,   2, 145,   1, 145,   0, 145,   0, 145,   0,  41,  31,  41,  30,  41,  29,  41,  28,  41,  27,  41,  26,  41,  25,  41,  24,  41,  23,  41,  22,  41,  21,  41,  20,  41,  19,  41,  18,  41,  17,  41,  16,  41,  15,  41,  14,  41,  13,  41,  12,  41,  11,  41,  10,  41,   9,  41,   8,  41,   7,  41,   6,  41,   5,  41,   4,  41,   3,  41,   2,  41,   1,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0, 244,  31, 244,  30, 244,  29, 244,  28, 244,  27, 244,  26, 244,  25, 244,  24, 218,  31, 218,  30, 218,  29, 218,  28, 218,  27, 218,  26, 218,  25, 218,  24, 218,  23, 218,  22, 218,  21, 218,  20, 218,  19, 218,  18, 218,  17, 218,  16, 218,  15, 218,  14, 218,  13, 218,  12, 218,  11, 218,  10, 218,   9, 218,   8, 218,   7, 218,   6, 218,   5, 218,   4, 218,   3, 218,   2, 218,   1, 218,   0, 218,   0, 218,   0, 218,   0, 218,   0, 218,   0, 218,   0, 218,   0, 218,   0, 218,   0, 218,   0, 218,   0, 218,   0, 218,   0, 218,   0, 218,   0, 218,   0, 218,   0, 144,  31, 144,  30, 144,  29, 144,  28, 144,  27, 144,  26, 144,  25, 144,  24, 144,  23, 144,  22, 144,  21, 144,  20, 144,  19, 144,  18, 144,  17, 144,  16, 144,  15, 144,  14, 144,  13, 144,  12, 144,  11, 144,  10, 144,   9, 144,   8, 144,   7, 144,   6, 144,   5, 144,   4, 144,   3, 144,   2, 144,   1, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0,  13,  31,  13,  30,  13,  29,  13,  28,  13,  27,  13,  26,  13,  25,  13,  24,  13,  23,  13,  22,  13,  21,  13,  20,  13,  19,  13,  18,  13,  17,  13,  16,  13,  15,  13,  14,  13,  13,  13,  12,  13,  11,  13,  10,  13,   9,  13,   8,  13,   7,  13,   6,  13,   5,  13,   4,  13,   3,  13,   2,  13,   1,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0, 160,  31, 160,  30, 160,  29, 160,  28, 160,  27, 160,  26, 160,  25, 160,  24, 160,  23, 160,  22, 160,  21, 160,  20, 160,  19, 160,  18, 160,  17, 160,  16, 160,  15, 160,  14, 160,  13, 160,  12, 160,  11, 160,  10, 160,   9, 160,   8, 160,   7, 160,   6, 160,   5, 160,   4, 160,   3, 160,   2, 160,   1, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 125,  31, 125,  30, 125,  29, 125,  28, 125,  27, 125,  26, 125,  25, 125,  24, 125,  23, 125,  22, 125,  21, 125,  20, 125,  19, 125,  18, 125,  17, 125,  16, 125,  15, 125,  14, 125,  13, 125,  12, 125,  11, 125,  10, 125,   9, 125,   8, 125,   7, 125,   6, 125,   5, 125,   4, 125,   3, 125,   2, 125,   1, 125,   0);
	constant SCENARIO_ADDRESS_1 : integer := 2056;


	--Scenario 2
	constant SCENARIO_LENGTH_2 : integer := 964;
	type scenario_type_2 is array (0 to SCENARIO_LENGTH_2*2-1) of integer;
	signal scenario_input_2 : scenario_type_2 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 222,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 244,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  15,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 179,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  75,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  66,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  28,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  55,   0,   0,   0, 151,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 170,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 194,   0,   0,   0, 215,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 207,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  13,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 249,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 106,   0, 246,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 213,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  86,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 147,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 194,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  84,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 120,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 184,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 127,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_2  : scenario_type_2 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 222,  31, 222,  30, 222,  29, 222,  28, 222,  27, 222,  26, 222,  25, 222,  24, 244,  31, 244,  30, 244,  29, 244,  28, 244,  27, 244,  26, 244,  25, 244,  24, 244,  23, 244,  22, 244,  21, 244,  20, 244,  19,  15,  31,  15,  30,  15,  29,  15,  28,  15,  27,  15,  26,  15,  25,  15,  24,  15,  23,  15,  22,  15,  21,  15,  20,  15,  19,  15,  18,  15,  17,  15,  16,  15,  15,  15,  14,  15,  13,  15,  12,  15,  11,  15,  10,  15,   9,  15,   8,  15,   7,  15,   6,  15,   5,  15,   4,  15,   3,  15,   2,  15,   1,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0, 179,  31, 179,  30, 179,  29, 179,  28, 179,  27, 179,  26, 179,  25, 179,  24, 179,  23, 179,  22, 179,  21, 179,  20, 179,  19, 179,  18, 179,  17, 179,  16, 179,  15, 179,  14, 179,  13, 179,  12, 179,  11, 179,  10, 179,   9, 179,   8, 179,   7, 179,   6, 179,   5, 179,   4, 179,   3, 179,   2, 179,   1,  75,  31,  75,  30,  75,  29,  75,  28,  75,  27,  75,  26,  75,  25,  75,  24,  75,  23,  75,  22,  75,  21,  75,  20,  75,  19,  75,  18,  75,  17,  75,  16,  75,  15,  75,  14,  75,  13,  75,  12,  75,  11,  75,  10,  66,  31,  66,  30,  66,  29,  66,  28,  66,  27,  66,  26,  66,  25,  66,  24,  66,  23,  66,  22,  66,  21,  66,  20,  66,  19,  66,  18,  66,  17,  66,  16,  66,  15,  66,  14,  66,  13,  66,  12,  66,  11,  66,  10,  66,   9,  66,   8,  66,   7,  66,   6,  66,   5,  66,   4,  66,   3,  66,   2,  66,   1,  66,   0,  66,   0,  66,   0,  66,   0,  66,   0,  66,   0,  66,   0,  66,   0,  66,   0,  66,   0,  66,   0,  66,   0,  66,   0,  66,   0,  66,   0,  66,   0,  66,   0,  66,   0,  66,   0,  28,  31,  28,  30,  28,  29,  28,  28,  28,  27,  28,  26,  28,  25,  28,  24,  28,  23,  28,  22,  28,  21,  28,  20,  28,  19,  28,  18,  28,  17,  28,  16,  28,  15,  28,  14,  28,  13,  28,  12,  28,  11,  28,  10,  28,   9,  28,   8,  28,   7,  28,   6,  28,   5,  28,   4,  28,   3,  28,   2,  28,   1,  28,   0,  28,   0,  28,   0,  28,   0,  28,   0,  28,   0,  28,   0,  28,   0,  28,   0,  28,   0,  28,   0,  28,   0,  28,   0,  28,   0,  28,   0,  55,  31,  55,  30, 151,  31, 151,  30, 151,  29, 151,  28, 151,  27, 151,  26, 151,  25, 151,  24, 151,  23, 151,  22, 151,  21, 151,  20, 151,  19, 151,  18, 151,  17, 151,  16, 151,  15, 151,  14, 151,  13, 151,  12, 151,  11, 151,  10, 151,   9, 151,   8, 151,   7, 170,  31, 170,  30, 170,  29, 170,  28, 170,  27, 170,  26, 170,  25, 170,  24, 170,  23, 170,  22, 170,  21, 170,  20, 170,  19, 170,  18, 170,  17, 170,  16, 170,  15, 170,  14, 170,  13, 194,  31, 194,  30, 215,  31, 215,  30, 215,  29, 215,  28, 215,  27, 215,  26, 215,  25, 215,  24, 215,  23, 215,  22, 215,  21, 215,  20, 215,  19, 215,  18, 215,  17, 215,  16, 215,  15, 215,  14, 215,  13, 215,  12, 215,  11, 215,  10, 215,   9, 215,   8, 215,   7, 215,   6, 215,   5, 215,   4, 215,   3, 215,   2, 215,   1, 215,   0, 215,   0, 215,   0, 215,   0, 215,   0, 215,   0, 215,   0, 215,   0, 215,   0, 215,   0, 215,   0, 215,   0, 215,   0, 215,   0, 215,   0, 215,   0, 215,   0, 215,   0, 215,   0, 215,   0, 215,   0, 215,   0, 215,   0, 215,   0, 207,  31, 207,  30, 207,  29, 207,  28, 207,  27, 207,  26, 207,  25, 207,  24, 207,  23, 207,  22, 207,  21, 207,  20, 207,  19, 207,  18, 207,  17, 207,  16, 207,  15, 207,  14, 207,  13, 207,  12, 207,  11, 207,  10,  13,  31,  13,  30,  13,  29,  13,  28,  13,  27,  13,  26,  13,  25,  13,  24,  13,  23,  13,  22,  13,  21,  13,  20,  13,  19,  13,  18,  13,  17,  13,  16,  13,  15,  13,  14,  13,  13,  13,  12,  13,  11,  13,  10,  13,   9,  13,   8, 249,  31, 249,  30, 249,  29, 249,  28, 249,  27, 249,  26, 249,  25, 249,  24, 249,  23, 249,  22, 249,  21, 249,  20, 249,  19, 249,  18, 106,  31, 246,  31, 246,  30, 246,  29, 246,  28, 246,  27, 246,  26, 246,  25, 246,  24, 246,  23, 246,  22, 246,  21, 246,  20, 246,  19, 246,  18, 246,  17, 246,  16, 246,  15, 246,  14, 246,  13, 246,  12, 246,  11, 213,  31, 213,  30, 213,  29, 213,  28, 213,  27, 213,  26, 213,  25, 213,  24, 213,  23, 213,  22,  86,  31,  86,  30,  86,  29,  86,  28,  86,  27,  86,  26,  86,  25,  86,  24,  86,  23,  86,  22,  86,  21,  86,  20,  86,  19,  86,  18,  86,  17,  86,  16,  86,  15,  86,  14,  86,  13,  86,  12,  86,  11,  86,  10,  86,   9,  86,   8,  86,   7,  86,   6,  86,   5,  86,   4,  86,   3,  86,   2,  86,   1,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0,  86,   0, 147,  31, 147,  30, 147,  29, 147,  28, 147,  27, 147,  26, 147,  25, 147,  24, 147,  23, 147,  22, 147,  21, 147,  20, 147,  19, 147,  18, 147,  17, 147,  16, 147,  15, 147,  14, 147,  13, 147,  12, 147,  11, 147,  10, 147,   9, 147,   8, 147,   7, 147,   6, 147,   5, 147,   4, 147,   3, 147,   2, 147,   1, 147,   0, 147,   0, 147,   0, 147,   0, 194,  31, 194,  30, 194,  29, 194,  28, 194,  27, 194,  26, 194,  25, 194,  24,  84,  31,  84,  30,  84,  29,  84,  28,  84,  27,  84,  26,  84,  25,  84,  24,  84,  23,  84,  22,  84,  21,  84,  20,  84,  19,  84,  18,  84,  17,  84,  16,  84,  15,  84,  14,  84,  13,  84,  12,  84,  11,  84,  10,  84,   9,  84,   8,  84,   7,  84,   6,  84,   5,  84,   4,  84,   3,  84,   2,  84,   1,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0,  84,   0, 120,  31, 120,  30, 120,  29, 120,  28, 120,  27, 120,  26, 120,  25, 120,  24, 120,  23, 120,  22, 120,  21, 120,  20, 120,  19, 120,  18, 120,  17, 120,  16, 120,  15, 120,  14, 120,  13, 120,  12, 120,  11, 120,  10, 120,   9, 120,   8, 120,   7, 120,   6, 120,   5, 120,   4, 120,   3, 120,   2, 120,   1, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 184,  31, 184,  30, 184,  29, 184,  28, 184,  27, 184,  26, 184,  25, 184,  24, 184,  23, 184,  22, 184,  21, 184,  20, 184,  19, 184,  18, 184,  17, 184,  16, 184,  15, 184,  14, 184,  13, 184,  12, 184,  11, 184,  10, 184,   9, 184,   8, 184,   7, 184,   6, 184,   5, 184,   4, 184,   3, 184,   2, 184,   1, 184,   0, 184,   0, 184,   0, 184,   0, 184,   0, 184,   0, 184,   0, 184,   0, 184,   0, 184,   0, 184,   0, 184,   0, 184,   0, 184,   0, 184,   0, 184,   0, 184,   0, 184,   0, 127,  31, 127,  30, 127,  29, 127,  28, 127,  27, 127,  26, 127,  25, 127,  24, 127,  23, 127,  22, 127,  21, 127,  20, 127,  19, 127,  18, 127,  17, 127,  16, 127,  15, 127,  14, 127,  13, 127,  12, 127,  11, 127,  10, 127,   9, 127,   8, 127,   7, 127,   6, 127,   5, 127,   4, 127,   3, 127,   2, 127,   1, 127,   0, 127,   0, 127,   0, 127,   0, 127,   0, 127,   0);
	constant SCENARIO_ADDRESS_2 : integer := 4154;


	--Scenario 3
	constant SCENARIO_LENGTH_3 : integer := 1023;
	type scenario_type_3 is array (0 to SCENARIO_LENGTH_3*2-1) of integer;
	signal scenario_input_3 : scenario_type_3 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 133,   0,   0,   0,   0,   0,  92,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 231,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 215,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 179,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 123,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 162,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  37,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 182,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  29,   0, 101,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 227,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 181,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 221,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  32,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  41,   0,  78,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 142,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  50,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 160,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 174,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 197,   0,   0,   0, 167,   0,   0,   0,   0,   0,   0,   0,   0,   0, 146,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 195,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  88,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  93,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  49,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 129,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  10,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  49,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 227,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 190,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  57,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_3  : scenario_type_3 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 133,  31, 133,  30, 133,  29,  92,  31,  92,  30,  92,  29,  92,  28,  92,  27,  92,  26,  92,  25,  92,  24,  92,  23,  92,  22,  92,  21,  92,  20,  92,  19,  92,  18,  92,  17,  92,  16,  92,  15,  92,  14,  92,  13,  92,  12,  92,  11,  92,  10,  92,   9,  92,   8, 231,  31, 231,  30, 231,  29, 231,  28, 231,  27, 231,  26, 231,  25, 231,  24, 215,  31, 215,  30, 215,  29, 215,  28, 215,  27, 215,  26, 215,  25, 179,  31, 179,  30, 179,  29, 179,  28, 179,  27, 179,  26, 179,  25, 179,  24, 179,  23, 179,  22, 179,  21, 179,  20, 179,  19, 179,  18, 179,  17, 179,  16, 179,  15, 179,  14, 179,  13, 179,  12, 179,  11, 179,  10, 179,   9, 179,   8, 179,   7, 179,   6, 179,   5, 179,   4, 179,   3, 179,   2, 179,   1, 123,  31, 123,  30, 123,  29, 123,  28, 123,  27, 123,  26, 123,  25, 123,  24, 123,  23, 123,  22, 123,  21, 123,  20, 123,  19, 123,  18, 123,  17, 123,  16, 123,  15, 123,  14, 123,  13, 123,  12, 123,  11, 123,  10, 123,   9, 123,   8, 123,   7, 123,   6, 123,   5, 123,   4, 123,   3, 123,   2, 123,   1, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 162,  31, 162,  30, 162,  29, 162,  28, 162,  27, 162,  26, 162,  25, 162,  24, 162,  23, 162,  22, 162,  21, 162,  20, 162,  19, 162,  18, 162,  17, 162,  16, 162,  15, 162,  14, 162,  13, 162,  12, 162,  11, 162,  10, 162,   9, 162,   8, 162,   7, 162,   6, 162,   5, 162,   4, 162,   3, 162,   2, 162,   1, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0,  37,  31,  37,  30,  37,  29,  37,  28,  37,  27,  37,  26,  37,  25,  37,  24,  37,  23,  37,  22,  37,  21,  37,  20,  37,  19,  37,  18,  37,  17,  37,  16,  37,  15,  37,  14,  37,  13,  37,  12,  37,  11,  37,  10,  37,   9,  37,   8,  37,   7,  37,   6,  37,   5,  37,   4,  37,   3,  37,   2,  37,   1,  37,   0,  37,   0,  37,   0,  37,   0,  37,   0,  37,   0,  37,   0,  37,   0, 182,  31, 182,  30, 182,  29, 182,  28, 182,  27, 182,  26, 182,  25, 182,  24, 182,  23, 182,  22, 182,  21, 182,  20, 182,  19, 182,  18, 182,  17, 182,  16, 182,  15, 182,  14, 182,  13, 182,  12, 182,  11, 182,  10, 182,   9, 182,   8, 182,   7, 182,   6, 182,   5, 182,   4, 182,   3, 182,   2, 182,   1, 182,   0, 182,   0, 182,   0, 182,   0, 182,   0, 182,   0, 182,   0, 182,   0, 182,   0, 182,   0, 182,   0, 182,   0, 182,   0, 182,   0, 182,   0, 182,   0, 182,   0, 182,   0,  29,  31, 101,  31, 101,  30, 101,  29, 101,  28, 101,  27, 101,  26, 101,  25, 101,  24, 101,  23, 101,  22, 101,  21, 101,  20, 101,  19, 101,  18, 101,  17, 101,  16, 101,  15, 101,  14, 101,  13, 101,  12, 101,  11, 101,  10, 101,   9, 101,   8, 101,   7, 101,   6, 101,   5, 101,   4, 101,   3, 101,   2, 101,   1, 101,   0, 101,   0, 101,   0, 101,   0, 101,   0, 101,   0, 101,   0, 101,   0, 101,   0, 101,   0, 101,   0, 101,   0, 101,   0, 101,   0, 101,   0, 101,   0, 101,   0, 101,   0, 101,   0, 101,   0, 101,   0, 101,   0, 101,   0, 227,  31, 227,  30, 227,  29, 227,  28, 227,  27, 227,  26, 227,  25, 227,  24, 227,  23, 227,  22, 227,  21, 227,  20, 227,  19, 227,  18, 227,  17, 227,  16, 227,  15, 227,  14, 227,  13, 227,  12, 227,  11, 227,  10, 227,   9, 227,   8, 227,   7, 227,   6, 227,   5, 227,   4, 227,   3, 227,   2, 227,   1, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 181,  31, 181,  30, 181,  29, 181,  28, 181,  27, 181,  26, 181,  25, 181,  24, 181,  23, 181,  22, 181,  21, 181,  20, 181,  19, 181,  18, 181,  17, 181,  16, 181,  15, 181,  14, 181,  13, 181,  12, 181,  11, 181,  10, 181,   9, 181,   8, 181,   7, 181,   6, 181,   5, 181,   4, 181,   3, 181,   2, 181,   1, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 181,   0, 221,  31, 221,  30, 221,  29, 221,  28, 221,  27, 221,  26, 221,  25, 221,  24, 221,  23, 221,  22, 221,  21,  32,  31,  32,  30,  32,  29,  32,  28,  32,  27,  32,  26,  32,  25,  32,  24,  32,  23,  32,  22,  32,  21,  32,  20,  32,  19,  32,  18,  32,  17,  32,  16,  32,  15,  32,  14,  32,  13,  32,  12,  32,  11,  32,  10,  32,   9,  32,   8,  32,   7,  32,   6,  32,   5,  32,   4,  32,   3,  32,   2,  32,   1,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  41,  31,  78,  31,  78,  30,  78,  29,  78,  28,  78,  27,  78,  26,  78,  25,  78,  24,  78,  23,  78,  22,  78,  21,  78,  20,  78,  19,  78,  18,  78,  17,  78,  16,  78,  15,  78,  14,  78,  13,  78,  12,  78,  11,  78,  10,  78,   9,  78,   8,  78,   7,  78,   6,  78,   5,  78,   4,  78,   3,  78,   2, 142,  31, 142,  30, 142,  29, 142,  28, 142,  27, 142,  26, 142,  25, 142,  24, 142,  23, 142,  22, 142,  21, 142,  20, 142,  19, 142,  18, 142,  17, 142,  16, 142,  15, 142,  14, 142,  13,  50,  31,  50,  30,  50,  29,  50,  28,  50,  27,  50,  26,  50,  25,  50,  24,  50,  23,  50,  22,  50,  21,  50,  20,  50,  19,  50,  18,  50,  17,  50,  16,  50,  15,  50,  14,  50,  13,  50,  12,  50,  11,  50,  10,  50,   9,  50,   8,  50,   7,  50,   6,  50,   5,  50,   4, 160,  31, 160,  30, 160,  29, 160,  28, 160,  27, 160,  26, 160,  25, 174,  31, 174,  30, 174,  29, 174,  28, 174,  27, 174,  26, 174,  25, 174,  24, 174,  23, 174,  22, 174,  21, 174,  20, 174,  19, 174,  18, 174,  17, 174,  16, 174,  15, 174,  14, 174,  13, 174,  12, 174,  11, 174,  10, 174,   9, 174,   8, 174,   7, 174,   6, 174,   5, 174,   4, 174,   3, 174,   2, 174,   1, 174,   0, 174,   0, 174,   0, 174,   0, 174,   0, 174,   0, 174,   0, 174,   0, 174,   0, 174,   0, 174,   0, 174,   0, 174,   0, 174,   0, 197,  31, 197,  30, 167,  31, 167,  30, 167,  29, 167,  28, 167,  27, 146,  31, 146,  30, 146,  29, 146,  28, 146,  27, 146,  26, 146,  25, 146,  24, 146,  23, 146,  22, 146,  21, 146,  20, 146,  19, 146,  18, 146,  17, 146,  16, 146,  15, 146,  14, 146,  13, 146,  12, 146,  11, 146,  10, 146,   9, 146,   8, 146,   7, 146,   6, 146,   5, 146,   4, 146,   3, 146,   2, 146,   1, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 195,  31, 195,  30, 195,  29, 195,  28, 195,  27, 195,  26, 195,  25,  88,  31,  88,  30,  88,  29,  88,  28,  88,  27,  88,  26,  88,  25,  88,  24,  88,  23,  88,  22,  88,  21,  88,  20,  88,  19,  88,  18,  88,  17,  88,  16,  88,  15,  88,  14,  88,  13,  88,  12,  88,  11,  88,  10,  88,   9,  88,   8,  88,   7,  88,   6,  88,   5,  88,   4,  88,   3,  88,   2,  88,   1,  88,   0,  88,   0,  88,   0,  93,  31,  93,  30,  93,  29,  93,  28,  93,  27,  93,  26,  93,  25,  93,  24,  49,  31,  49,  30,  49,  29,  49,  28,  49,  27,  49,  26,  49,  25,  49,  24,  49,  23,  49,  22,  49,  21,  49,  20,  49,  19,  49,  18,  49,  17,  49,  16,  49,  15,  49,  14,  49,  13,  49,  12,  49,  11,  49,  10,  49,   9,  49,   8,  49,   7,  49,   6,  49,   5,  49,   4,  49,   3, 129,  31, 129,  30, 129,  29, 129,  28, 129,  27, 129,  26, 129,  25, 129,  24, 129,  23, 129,  22, 129,  21, 129,  20, 129,  19, 129,  18, 129,  17, 129,  16, 129,  15, 129,  14, 129,  13, 129,  12, 129,  11, 129,  10, 129,   9, 129,   8, 129,   7, 129,   6, 129,   5,  10,  31,  10,  30,  10,  29,  10,  28,  10,  27,  10,  26,  10,  25,  10,  24,  10,  23,  10,  22,  10,  21,  10,  20,  10,  19,  10,  18,  10,  17,  10,  16,  10,  15,  10,  14,  10,  13,  10,  12,  10,  11,  10,  10,  10,   9,  10,   8,  10,   7,  10,   6,  10,   5,  10,   4,  10,   3,  10,   2,  10,   1,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  49,  31,  49,  30,  49,  29,  49,  28,  49,  27,  49,  26,  49,  25,  49,  24,  49,  23,  49,  22,  49,  21,  49,  20,  49,  19,  49,  18,  49,  17,  49,  16,  49,  15,  49,  14,  49,  13,  49,  12,  49,  11,  49,  10,  49,   9,  49,   8,  49,   7,  49,   6,  49,   5,  49,   4,  49,   3,  49,   2,  49,   1,  49,   0,  49,   0,  49,   0,  49,   0,  49,   0,  49,   0,  49,   0,  49,   0,  49,   0,  49,   0,  49,   0,  49,   0,  49,   0,  49,   0,  49,   0,  49,   0,  49,   0, 227,  31, 227,  30, 227,  29, 227,  28, 227,  27, 227,  26, 227,  25, 227,  24, 227,  23, 227,  22, 227,  21, 227,  20, 227,  19, 227,  18, 227,  17, 227,  16, 227,  15, 227,  14, 227,  13, 227,  12, 227,  11, 227,  10, 227,   9, 227,   8, 227,   7, 227,   6, 227,   5, 227,   4, 227,   3, 227,   2, 227,   1, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 190,  31, 190,  30, 190,  29, 190,  28, 190,  27, 190,  26, 190,  25, 190,  24,  57,  31,  57,  30,  57,  29,  57,  28,  57,  27,  57,  26,  57,  25,  57,  24,  57,  23,  57,  22,  57,  21,  57,  20,  57,  19,  57,  18,  57,  17,  57,  16,  57,  15,  57,  14,  57,  13,  57,  12,  57,  11,  57,  10,  57,   9,  57,   8,  57,   7,  57,   6,  57,   5,  57,   4,  57,   3,  57,   2,  57,   1,  57,   0,  57,   0,  57,   0,  57,   0,  57,   0,  57,   0,  57,   0,  57,   0,  57,   0,  57,   0,  57,   0,  57,   0);
	constant SCENARIO_ADDRESS_3 : integer := 6145;


	--Scenario 4
	constant SCENARIO_LENGTH_4 : integer := 1;
	type scenario_type_4 is array (0 to SCENARIO_LENGTH_4*2-1) of integer;
	signal scenario_input_4 : scenario_type_4 := (7,   7);
	signal scenario_full_4  : scenario_type_4 := (7,   7);
	constant SCENARIO_ADDRESS_4 : integer := 10099;
	--This sequence is going to be ignored by the component
	--as the i_k parameter is will be set to zero


	--Scenario 5
	constant SCENARIO_LENGTH_5 : integer := 1021;
	type scenario_type_5 is array (0 to SCENARIO_LENGTH_5*2-1) of integer;
	signal scenario_input_5 : scenario_type_5 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  58,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 180,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 122,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 204,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  65,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  32,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  18,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 121,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  81,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 179,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  78,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  27,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 146,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 130,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  89,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  62,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  72,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  93,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 126,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 243,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 114,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 246,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  14,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  32,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 142,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_5  : scenario_type_5 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  58,  31,  58,  30,  58,  29,  58,  28,  58,  27,  58,  26,  58,  25,  58,  24,  58,  23,  58,  22,  58,  21,  58,  20,  58,  19,  58,  18,  58,  17,  58,  16,  58,  15,  58,  14,  58,  13,  58,  12,  58,  11,  58,  10,  58,   9,  58,   8,  58,   7,  58,   6,  58,   5,  58,   4,  58,   3, 180,  31, 180,  30, 180,  29, 180,  28, 180,  27, 180,  26, 180,  25, 180,  24, 180,  23, 180,  22, 180,  21, 180,  20, 180,  19, 180,  18, 180,  17, 180,  16, 180,  15, 180,  14, 180,  13, 180,  12, 180,  11, 180,  10, 180,   9, 180,   8, 180,   7, 180,   6, 180,   5, 180,   4, 180,   3, 180,   2, 180,   1, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 122,  31, 122,  30, 122,  29, 122,  28, 122,  27, 122,  26, 122,  25, 122,  24, 122,  23, 122,  22, 122,  21, 122,  20, 122,  19, 122,  18, 122,  17, 122,  16, 122,  15, 122,  14, 122,  13, 204,  31, 204,  30, 204,  29, 204,  28, 204,  27, 204,  26, 204,  25, 204,  24, 204,  23, 204,  22, 204,  21, 204,  20, 204,  19, 204,  18, 204,  17, 204,  16, 204,  15, 204,  14, 204,  13, 204,  12, 204,  11, 204,  10, 204,   9, 204,   8, 204,   7, 204,   6, 204,   5, 204,   4, 204,   3, 204,   2, 204,   1, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0,  65,  31,  65,  30,  65,  29,  65,  28,  65,  27,  65,  26,  65,  25,  65,  24,  65,  23,  65,  22,  65,  21,  65,  20,  65,  19,  65,  18,  65,  17,  65,  16,  65,  15,  65,  14,  65,  13,  65,  12,  65,  11,  65,  10,  65,   9,  65,   8,  65,   7,  65,   6,  65,   5,  65,   4,  65,   3,  65,   2,  65,   1,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  32,  31,  32,  30,  32,  29,  32,  28,  32,  27,  32,  26,  32,  25,  32,  24,  32,  23,  32,  22,  32,  21,  32,  20,  32,  19,  32,  18,  32,  17,  32,  16,  32,  15,  32,  14,  32,  13,  32,  12,  32,  11,  32,  10,  32,   9,  32,   8,  18,  31,  18,  30,  18,  29,  18,  28,  18,  27,  18,  26, 121,  31, 121,  30, 121,  29, 121,  28, 121,  27, 121,  26, 121,  25, 121,  24, 121,  23, 121,  22, 121,  21, 121,  20, 121,  19, 121,  18, 121,  17, 121,  16, 121,  15, 121,  14, 121,  13, 121,  12, 121,  11, 121,  10, 121,   9, 121,   8, 121,   7, 121,   6, 121,   5, 121,   4, 121,   3, 121,   2, 121,   1, 121,   0, 121,   0, 121,   0, 121,   0,  81,  31,  81,  30,  81,  29,  81,  28,  81,  27,  81,  26,  81,  25,  81,  24,  81,  23,  81,  22,  81,  21,  81,  20,  81,  19,  81,  18,  81,  17,  81,  16,  81,  15,  81,  14,  81,  13,  81,  12,  81,  11,  81,  10,  81,   9,  81,   8,  81,   7, 179,  31, 179,  30, 179,  29, 179,  28, 179,  27, 179,  26, 179,  25, 179,  24, 179,  23, 179,  22, 179,  21, 179,  20, 179,  19, 179,  18, 179,  17, 179,  16, 179,  15, 179,  14, 179,  13, 179,  12, 179,  11, 179,  10, 179,   9, 179,   8, 179,   7, 179,   6, 179,   5, 179,   4, 179,   3, 179,   2, 179,   1, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0,  78,  31,  78,  30,  78,  29,  78,  28,  78,  27,  78,  26,  78,  25,  78,  24,  78,  23,  78,  22,  78,  21,  78,  20,  78,  19,  78,  18,  78,  17,  78,  16,  78,  15,  78,  14,  78,  13,  78,  12,  78,  11,  78,  10,  78,   9,  78,   8,  78,   7,  78,   6,  78,   5,  78,   4,  78,   3,  78,   2,  78,   1,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  27,  31,  27,  30,  27,  29,  27,  28,  27,  27,  27,  26,  27,  25,  27,  24,  27,  23,  27,  22, 146,  31, 146,  30, 146,  29, 146,  28, 146,  27, 146,  26, 146,  25, 146,  24, 146,  23, 146,  22, 146,  21, 146,  20, 146,  19, 146,  18, 146,  17, 146,  16, 146,  15, 146,  14, 146,  13, 146,  12, 146,  11, 146,  10, 146,   9, 146,   8, 146,   7, 146,   6, 146,   5, 146,   4, 146,   3, 146,   2, 146,   1, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 130,  31, 130,  30, 130,  29, 130,  28, 130,  27, 130,  26, 130,  25, 130,  24, 130,  23, 130,  22, 130,  21, 130,  20, 130,  19, 130,  18, 130,  17, 130,  16, 130,  15, 130,  14, 130,  13, 130,  12, 130,  11, 130,  10, 130,   9, 130,   8, 130,   7, 130,   6, 130,   5, 130,   4, 130,   3, 130,   2, 130,   1, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0,  89,  31,  89,  30,  89,  29,  89,  28,  89,  27,  89,  26,  89,  25,  89,  24,  89,  23,  89,  22,  62,  31,  62,  30,  62,  29,  62,  28,  62,  27,  62,  26,  62,  25,  62,  24,  62,  23,  62,  22,  62,  21,  62,  20,  62,  19,  62,  18,  62,  17,  62,  16,  62,  15,  62,  14,  62,  13,  62,  12,  62,  11,  62,  10,  62,   9,  62,   8,  62,   7,  62,   6,  62,   5,  62,   4,  62,   3,  62,   2,  62,   1,  72,  31,  72,  30,  72,  29,  72,  28,  72,  27,  72,  26,  72,  25,  72,  24,  72,  23,  72,  22,  72,  21,  72,  20,  72,  19,  72,  18,  72,  17,  72,  16,  72,  15,  72,  14,  72,  13,  72,  12,  72,  11,  72,  10,  72,   9,  72,   8,  93,  31,  93,  30,  93,  29,  93,  28,  93,  27,  93,  26,  93,  25,  93,  24,  93,  23,  93,  22,  93,  21,  93,  20,  93,  19,  93,  18,  93,  17,  93,  16,  93,  15,  93,  14,  93,  13,  93,  12,  93,  11,  93,  10,  93,   9,  93,   8,  93,   7,  93,   6,  93,   5,  93,   4,  93,   3,  93,   2,  93,   1, 126,  31, 126,  30, 126,  29, 126,  28, 126,  27, 126,  26, 126,  25, 126,  24, 126,  23, 126,  22, 126,  21, 126,  20, 126,  19, 126,  18, 126,  17, 126,  16, 126,  15, 126,  14, 126,  13, 126,  12, 126,  11, 126,  10, 126,   9, 126,   8, 126,   7, 126,   6, 126,   5, 126,   4, 126,   3, 126,   2, 126,   1, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 126,   0, 243,  31, 243,  30, 243,  29, 243,  28, 243,  27, 243,  26, 243,  25, 243,  24, 243,  23, 243,  22, 243,  21, 243,  20, 243,  19, 243,  18, 243,  17, 243,  16, 243,  15, 243,  14, 243,  13, 243,  12, 243,  11, 243,  10, 243,   9, 243,   8, 243,   7, 243,   6, 243,   5, 243,   4, 243,   3, 243,   2, 114,  31, 114,  30, 114,  29, 114,  28, 114,  27, 114,  26, 114,  25, 114,  24, 114,  23, 114,  22, 114,  21, 114,  20, 114,  19, 114,  18, 114,  17, 114,  16, 114,  15, 114,  14, 114,  13, 114,  12, 114,  11, 114,  10, 114,   9, 114,   8, 114,   7, 114,   6, 114,   5, 246,  31, 246,  30, 246,  29, 246,  28, 246,  27, 246,  26, 246,  25, 246,  24, 246,  23, 246,  22, 246,  21, 246,  20, 246,  19, 246,  18, 246,  17, 246,  16, 246,  15, 246,  14, 246,  13, 246,  12, 246,  11, 246,  10, 246,   9, 246,   8, 246,   7, 246,   6, 246,   5, 246,   4, 246,   3, 246,   2, 246,   1, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0,  14,  31,  14,  30,  14,  29,  14,  28,  14,  27,  14,  26,  14,  25,  14,  24,  14,  23,  14,  22,  14,  21,  14,  20,  14,  19,  14,  18,  14,  17,  14,  16,  14,  15,  32,  31,  32,  30,  32,  29,  32,  28,  32,  27,  32,  26,  32,  25,  32,  24,  32,  23,  32,  22,  32,  21,  32,  20,  32,  19,  32,  18,  32,  17,  32,  16,  32,  15,  32,  14, 142,  31, 142,  30, 142,  29, 142,  28, 142,  27, 142,  26, 142,  25, 142,  24, 142,  23, 142,  22, 142,  21, 142,  20, 142,  19, 142,  18, 142,  17, 142,  16, 142,  15, 142,  14, 142,  13, 142,  12, 142,  11, 142,  10, 142,   9, 142,   8, 142,   7, 142,   6, 142,   5, 142,   4, 142,   3, 142,   2, 142,   1, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0);
	constant SCENARIO_ADDRESS_5 : integer := 10240;


	--Scenario 6
	constant SCENARIO_LENGTH_6 : integer := 983;
	type scenario_type_6 is array (0 to SCENARIO_LENGTH_6*2-1) of integer;
	signal scenario_input_6 : scenario_type_6 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 110,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 238,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 245,   0,   0,   0,   0,   0,  18,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 195,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 218,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 171,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 147,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  82,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 195,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 152,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  56,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 128,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 182,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  84,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 162,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 144,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 171,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 217,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  77,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  62,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  63,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 131,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 150,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 178,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  19,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 192,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_6  : scenario_type_6 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 110,  31, 110,  30, 110,  29, 110,  28, 110,  27, 110,  26, 110,  25, 110,  24, 110,  23, 110,  22, 110,  21, 110,  20, 110,  19, 110,  18, 110,  17, 110,  16, 110,  15, 110,  14, 110,  13, 110,  12, 110,  11, 110,  10, 110,   9, 110,   8, 110,   7, 110,   6, 110,   5, 110,   4, 110,   3, 110,   2, 110,   1, 110,   0, 110,   0, 110,   0, 110,   0, 110,   0, 110,   0, 110,   0, 110,   0, 110,   0, 110,   0, 110,   0, 110,   0, 110,   0, 110,   0, 110,   0, 110,   0, 110,   0, 110,   0, 238,  31, 238,  30, 238,  29, 238,  28, 238,  27, 238,  26, 238,  25, 238,  24, 238,  23, 238,  22, 245,  31, 245,  30, 245,  29,  18,  31,  18,  30,  18,  29,  18,  28,  18,  27,  18,  26,  18,  25,  18,  24,  18,  23,  18,  22,  18,  21,  18,  20,  18,  19,  18,  18,  18,  17,  18,  16,  18,  15,  18,  14,  18,  13,  18,  12,  18,  11,  18,  10,  18,   9,  18,   8, 195,  31, 195,  30, 195,  29, 195,  28, 195,  27, 195,  26, 195,  25, 195,  24, 195,  23, 195,  22, 195,  21, 195,  20, 195,  19, 195,  18, 195,  17, 195,  16, 195,  15, 195,  14, 195,  13, 195,  12, 195,  11, 195,  10, 195,   9, 195,   8, 195,   7, 195,   6, 195,   5, 195,   4, 195,   3, 195,   2, 195,   1, 195,   0, 195,   0, 195,   0, 195,   0, 195,   0, 195,   0, 195,   0, 195,   0, 195,   0, 195,   0, 195,   0, 195,   0, 195,   0, 195,   0, 195,   0, 218,  31, 218,  30, 218,  29, 218,  28, 218,  27, 218,  26, 218,  25, 218,  24, 218,  23, 218,  22, 171,  31, 171,  30, 171,  29, 171,  28, 171,  27, 171,  26, 171,  25, 171,  24, 171,  23, 171,  22, 171,  21, 171,  20, 171,  19, 171,  18, 171,  17, 171,  16, 171,  15, 171,  14, 171,  13, 171,  12, 171,  11, 171,  10, 171,   9, 147,  31, 147,  30, 147,  29, 147,  28, 147,  27, 147,  26, 147,  25, 147,  24, 147,  23, 147,  22, 147,  21, 147,  20, 147,  19, 147,  18, 147,  17, 147,  16, 147,  15, 147,  14, 147,  13, 147,  12, 147,  11, 147,  10, 147,   9, 147,   8, 147,   7, 147,   6, 147,   5, 147,   4, 147,   3, 147,   2, 147,   1, 147,   0, 147,   0, 147,   0,  82,  31,  82,  30,  82,  29,  82,  28,  82,  27,  82,  26,  82,  25,  82,  24,  82,  23,  82,  22,  82,  21,  82,  20,  82,  19,  82,  18,  82,  17,  82,  16,  82,  15,  82,  14, 195,  31, 195,  30, 195,  29, 195,  28, 195,  27, 195,  26, 195,  25, 195,  24, 152,  31, 152,  30, 152,  29, 152,  28, 152,  27, 152,  26, 152,  25, 152,  24, 152,  23, 152,  22, 152,  21, 152,  20, 152,  19, 152,  18, 152,  17, 152,  16, 152,  15, 152,  14, 152,  13, 152,  12, 152,  11, 152,  10, 152,   9, 152,   8, 152,   7, 152,   6, 152,   5, 152,   4, 152,   3, 152,   2, 152,   1, 152,   0, 152,   0, 152,   0, 152,   0, 152,   0, 152,   0, 152,   0, 152,   0,  56,  31,  56,  30,  56,  29,  56,  28,  56,  27,  56,  26,  56,  25,  56,  24,  56,  23,  56,  22,  56,  21,  56,  20,  56,  19,  56,  18,  56,  17,  56,  16,  56,  15,  56,  14,  56,  13,  56,  12,  56,  11,  56,  10,  56,   9,  56,   8,  56,   7,  56,   6,  56,   5, 128,  31, 128,  30, 128,  29, 128,  28, 128,  27, 128,  26, 128,  25, 128,  24, 128,  23, 128,  22, 128,  21, 128,  20, 128,  19, 128,  18, 128,  17, 128,  16, 128,  15, 128,  14, 128,  13, 128,  12, 128,  11, 128,  10, 128,   9, 128,   8, 128,   7, 128,   6, 128,   5, 128,   4, 128,   3, 128,   2, 128,   1, 128,   0, 128,   0, 128,   0, 128,   0, 128,   0, 128,   0, 128,   0, 182,  31, 182,  30, 182,  29, 182,  28, 182,  27, 182,  26, 182,  25, 182,  24, 182,  23, 182,  22, 182,  21, 182,  20, 182,  19, 182,  18, 182,  17, 182,  16, 182,  15, 182,  14, 182,  13, 182,  12, 182,  11, 182,  10, 182,   9, 182,   8, 182,   7, 182,   6, 182,   5, 182,   4, 182,   3, 182,   2, 182,   1,  84,  31,  84,  30,  84,  29,  84,  28,  84,  27,  84,  26,  84,  25,  84,  24,  84,  23,  84,  22,  84,  21,  84,  20,  84,  19,  84,  18,  84,  17,  84,  16,  84,  15,  84,  14,  84,  13,  84,  12, 162,  31, 162,  30, 162,  29, 162,  28, 162,  27, 162,  26, 162,  25, 162,  24, 162,  23, 162,  22, 162,  21, 162,  20, 162,  19, 162,  18, 162,  17, 162,  16, 162,  15, 162,  14, 162,  13, 162,  12, 162,  11, 162,  10, 162,   9, 162,   8, 162,   7, 162,   6, 162,   5, 162,   4, 162,   3, 162,   2, 162,   1, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 144,  31, 144,  30, 144,  29, 144,  28, 144,  27, 144,  26, 144,  25, 144,  24, 144,  23, 144,  22, 144,  21, 144,  20, 144,  19, 144,  18, 144,  17, 144,  16, 144,  15, 144,  14, 144,  13, 144,  12, 144,  11, 144,  10, 144,   9, 144,   8, 144,   7, 144,   6, 144,   5, 144,   4, 144,   3, 144,   2, 144,   1, 144,   0, 171,  31, 171,  30, 171,  29, 171,  28, 171,  27, 171,  26, 171,  25, 171,  24, 171,  23, 171,  22, 171,  21, 171,  20, 171,  19, 171,  18, 171,  17, 171,  16, 171,  15, 171,  14, 171,  13, 171,  12, 171,  11, 171,  10, 171,   9, 171,   8, 171,   7, 171,   6, 171,   5, 217,  31, 217,  30, 217,  29, 217,  28, 217,  27, 217,  26, 217,  25, 217,  24, 217,  23, 217,  22, 217,  21, 217,  20, 217,  19, 217,  18, 217,  17, 217,  16, 217,  15, 217,  14, 217,  13,  77,  31,  77,  30,  77,  29,  77,  28,  77,  27,  77,  26,  77,  25,  77,  24,  77,  23,  77,  22,  77,  21,  77,  20,  77,  19,  77,  18,  77,  17,  77,  16,  77,  15,  77,  14,  77,  13,  77,  12,  77,  11,  77,  10,  77,   9,  77,   8,  77,   7,  77,   6,  77,   5,  77,   4,  77,   3,  77,   2,  77,   1,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  77,   0,  62,  31,  62,  30,  62,  29,  62,  28,  62,  27,  62,  26,  62,  25,  62,  24,  62,  23,  62,  22,  62,  21,  62,  20,  62,  19,  62,  18,  62,  17,  62,  16,  62,  15,  62,  14,  62,  13,  62,  12,  62,  11,  62,  10,  62,   9,  62,   8,  62,   7,  62,   6,  62,   5,  62,   4,  62,   3,  62,   2,  62,   1,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  63,  31,  63,  30,  63,  29,  63,  28,  63,  27,  63,  26,  63,  25,  63,  24,  63,  23,  63,  22,  63,  21,  63,  20, 131,  31, 131,  30, 131,  29, 131,  28, 131,  27, 131,  26, 131,  25, 131,  24, 131,  23, 131,  22, 131,  21, 131,  20, 131,  19, 131,  18, 131,  17, 131,  16, 131,  15, 131,  14, 131,  13, 131,  12, 131,  11, 131,  10, 131,   9, 131,   8, 131,   7, 131,   6, 131,   5, 131,   4, 131,   3, 131,   2, 131,   1, 131,   0, 131,   0, 131,   0, 131,   0, 131,   0, 150,  31, 150,  30, 150,  29, 150,  28, 150,  27, 150,  26, 150,  25, 150,  24, 150,  23, 150,  22, 150,  21, 150,  20, 150,  19, 150,  18, 150,  17, 150,  16, 150,  15, 150,  14, 150,  13, 150,  12, 150,  11, 150,  10, 150,   9, 150,   8, 150,   7, 150,   6, 150,   5, 150,   4, 150,   3, 150,   2, 150,   1, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 178,  31, 178,  30, 178,  29, 178,  28, 178,  27, 178,  26, 178,  25, 178,  24, 178,  23,  19,  31,  19,  30,  19,  29,  19,  28,  19,  27,  19,  26,  19,  25,  19,  24,  19,  23,  19,  22,  19,  21,  19,  20,  19,  19,  19,  18,  19,  17,  19,  16,  19,  15,  19,  14,  19,  13,  19,  12,  19,  11,  19,  10,  19,   9, 192,  31, 192,  30, 192,  29, 192,  28, 192,  27, 192,  26, 192,  25, 192,  24, 192,  23, 192,  22, 192,  21, 192,  20, 192,  19, 192,  18, 192,  17, 192,  16, 192,  15, 192,  14, 192,  13, 192,  12, 192,  11, 192,  10, 192,   9, 192,   8, 192,   7, 192,   6, 192,   5, 192,   4, 192,   3, 192,   2, 192,   1, 192,   0, 192,   0, 192,   0, 192,   0, 192,   0, 192,   0, 192,   0, 192,   0, 192,   0, 192,   0, 192,   0, 192,   0, 192,   0, 192,   0, 192,   0, 192,   0, 192,   0, 192,   0, 192,   0, 192,   0, 192,   0);
	constant SCENARIO_ADDRESS_6 : integer := 12324;


	--Scenario 7
	constant SCENARIO_LENGTH_7 : integer := 1016;
	type scenario_type_7 is array (0 to SCENARIO_LENGTH_7*2-1) of integer;
	signal scenario_input_7 : scenario_type_7 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 212,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 190,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  64,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  58,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 197,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 127,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 183,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 100,   0,   0,   0, 100,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 214,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 194,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 239,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 204,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  55,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 106,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 210,   0,   0,   0,  95,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 125,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  35,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  26,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  11,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_7  : scenario_type_7 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 212,  31, 212,  30, 212,  29, 212,  28, 212,  27, 212,  26, 212,  25, 212,  24, 212,  23, 212,  22, 212,  21, 212,  20, 212,  19, 212,  18, 212,  17, 212,  16, 212,  15, 212,  14, 212,  13, 212,  12, 212,  11, 212,  10, 190,  31, 190,  30, 190,  29, 190,  28, 190,  27, 190,  26, 190,  25, 190,  24, 190,  23, 190,  22, 190,  21, 190,  20, 190,  19, 190,  18, 190,  17, 190,  16, 190,  15, 190,  14, 190,  13, 190,  12, 190,  11, 190,  10, 190,   9, 190,   8, 190,   7, 190,   6, 190,   5, 190,   4, 190,   3, 190,   2, 190,   1, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0,  64,  31,  64,  30,  64,  29,  64,  28,  64,  27,  64,  26,  64,  25,  64,  24,  64,  23,  64,  22,  64,  21,  64,  20,  64,  19,  64,  18,  64,  17,  64,  16,  64,  15,  64,  14,  64,  13,  64,  12,  64,  11,  64,  10,  64,   9,  64,   8,  64,   7,  64,   6,  64,   5,  64,   4,  64,   3,  64,   2,  64,   1,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  58,  31,  58,  30,  58,  29,  58,  28,  58,  27,  58,  26,  58,  25,  58,  24,  58,  23,  58,  22,  58,  21,  58,  20,  58,  19,  58,  18,  58,  17,  58,  16,  58,  15,  58,  14,  58,  13,  58,  12,  58,  11,  58,  10,  58,   9,  58,   8,  58,   7,  58,   6,  58,   5,  58,   4,  58,   3, 197,  31, 197,  30, 197,  29, 197,  28, 197,  27, 197,  26, 197,  25, 197,  24, 197,  23, 197,  22, 197,  21, 197,  20, 197,  19, 197,  18, 197,  17, 197,  16, 197,  15, 197,  14, 197,  13, 197,  12, 197,  11, 197,  10, 197,   9, 197,   8, 197,   7, 197,   6, 197,   5, 197,   4, 197,   3, 197,   2, 197,   1, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 127,  31, 127,  30, 127,  29, 127,  28, 127,  27, 127,  26, 127,  25, 127,  24, 127,  23, 127,  22, 127,  21, 127,  20, 127,  19, 127,  18, 127,  17, 127,  16, 127,  15, 127,  14, 127,  13, 127,  12, 127,  11, 127,  10, 127,   9, 127,   8, 127,   7, 127,   6, 127,   5, 127,   4, 127,   3, 127,   2, 183,  31, 183,  30, 183,  29, 183,  28, 183,  27, 183,  26, 183,  25, 183,  24, 183,  23, 183,  22, 183,  21, 183,  20, 183,  19, 183,  18, 183,  17, 183,  16, 183,  15, 183,  14, 183,  13, 183,  12, 183,  11, 183,  10, 183,   9, 183,   8, 183,   7, 183,   6, 183,   5, 183,   4, 183,   3, 183,   2, 183,   1, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 100,  31, 100,  30, 100,  31, 100,  30, 100,  29, 100,  28, 100,  27, 100,  26, 100,  25, 100,  24, 100,  23, 100,  22, 100,  21, 100,  20, 100,  19, 100,  18, 100,  17, 100,  16, 100,  15, 100,  14, 100,  13, 100,  12, 100,  11, 100,  10, 100,   9, 100,   8, 100,   7, 100,   6, 214,  31, 214,  30, 214,  29, 214,  28, 214,  27, 214,  26, 214,  25, 214,  24, 214,  23, 214,  22, 214,  21, 214,  20, 214,  19, 214,  18, 214,  17, 214,  16, 214,  15, 214,  14, 214,  13, 214,  12, 214,  11, 214,  10, 214,   9, 214,   8, 214,   7, 214,   6, 214,   5, 214,   4, 214,   3, 214,   2, 214,   1, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 194,  31, 194,  30, 194,  29, 194,  28, 194,  27, 194,  26, 194,  25, 194,  24, 194,  23, 194,  22, 194,  21, 194,  20, 194,  19, 194,  18, 194,  17, 194,  16, 194,  15, 194,  14, 194,  13, 194,  12, 194,  11, 194,  10, 194,   9, 194,   8, 194,   7, 194,   6, 194,   5, 194,   4, 194,   3, 194,   2, 194,   1, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 239,  31, 239,  30, 239,  29, 239,  28, 239,  27, 239,  26, 239,  25, 239,  24, 239,  23, 239,  22, 239,  21, 239,  20, 239,  19, 239,  18, 239,  17, 239,  16, 239,  15, 239,  14, 239,  13, 239,  12, 239,  11, 239,  10, 239,   9, 239,   8, 239,   7, 239,   6, 239,   5, 239,   4, 239,   3, 204,  31, 204,  30, 204,  29, 204,  28, 204,  27, 204,  26, 204,  25, 204,  24, 204,  23, 204,  22, 204,  21, 204,  20, 204,  19, 204,  18, 204,  17, 204,  16, 204,  15, 204,  14, 204,  13, 204,  12, 204,  11, 204,  10, 204,   9, 204,   8, 204,   7, 204,   6, 204,   5, 204,   4, 204,   3,  55,  31,  55,  30,  55,  29,  55,  28,  55,  27,  55,  26,  55,  25,  55,  24,  55,  23,  55,  22,  55,  21,  55,  20,  55,  19,  55,  18,  55,  17,  55,  16,  55,  15,  55,  14,  55,  13,  55,  12,  55,  11,  55,  10, 106,  31, 106,  30, 106,  29, 106,  28, 106,  27, 106,  26, 106,  25, 106,  24, 106,  23, 106,  22, 106,  21, 106,  20, 106,  19, 106,  18, 106,  17, 106,  16, 106,  15, 106,  14, 106,  13, 106,  12, 106,  11, 106,  10, 106,   9, 106,   8, 106,   7, 106,   6, 106,   5, 106,   4, 106,   3, 106,   2, 106,   1, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 106,   0, 210,  31, 210,  30,  95,  31,  95,  30,  95,  29,  95,  28,  95,  27,  95,  26,  95,  25,  95,  24,  95,  23,  95,  22,  95,  21,  95,  20,  95,  19,  95,  18,  95,  17,  95,  16,  95,  15,  95,  14,  95,  13,  95,  12,  95,  11,  95,  10,  95,   9,  95,   8,  95,   7,  95,   6,  95,   5,  95,   4,  95,   3,  95,   2, 125,  31, 125,  30, 125,  29, 125,  28, 125,  27, 125,  26, 125,  25, 125,  24, 125,  23, 125,  22, 125,  21, 125,  20, 125,  19, 125,  18, 125,  17, 125,  16, 125,  15, 125,  14, 125,  13, 125,  12, 125,  11, 125,  10, 125,   9, 125,   8, 125,   7, 125,   6, 125,   5,  35,  31,  35,  30,  35,  29,  35,  28,  35,  27,  35,  26,  35,  25,  35,  24,  35,  23,  35,  22,  35,  21,  35,  20,  26,  31,  26,  30,  26,  29,  26,  28,  26,  27,  26,  26,  26,  25,  26,  24,  26,  23,  26,  22,  26,  21,  26,  20,  26,  19,  26,  18,  26,  17,  26,  16,  26,  15,  26,  14,  26,  13,  26,  12,  26,  11,  26,  10,  26,   9,  26,   8,  26,   7,  26,   6,  26,   5,  26,   4,  26,   3,  26,   2,  26,   1,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  26,   0,  11,  31,  11,  30,  11,  29,  11,  28,  11,  27,  11,  26,  11,  25,  11,  24,  11,  23,  11,  22,  11,  21,  11,  20,  11,  19,  11,  18,  11,  17,  11,  16,  11,  15,  11,  14,  11,  13,  11,  12,  11,  11,  11,  10,  11,   9,  11,   8,  11,   7,  11,   6,  11,   5,  11,   4,  11,   3,  11,   2,  11,   1,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0);
	constant SCENARIO_ADDRESS_7 : integer := 14342;


	--Scenario 8
	constant SCENARIO_LENGTH_8 : integer := 1;
	type scenario_type_8 is array (0 to SCENARIO_LENGTH_8*2-1) of integer;
	signal scenario_input_8 : scenario_type_8 := (7,   7);
	signal scenario_full_8  : scenario_type_8 := (7,   7);
	constant SCENARIO_ADDRESS_8 : integer := 17055;
	--This sequence is going to be ignored by the component
	--as the i_k parameter is will be set to zero


	--Scenario 9
	constant SCENARIO_LENGTH_9 : integer := 1016;
	type scenario_type_9 is array (0 to SCENARIO_LENGTH_9*2-1) of integer;
	signal scenario_input_9 : scenario_type_9 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  31,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 230,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  33,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  21,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  87,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 200,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  58,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 152,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 129,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 228,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   6,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 250,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 179,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 151,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 241,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 133,   0,   0,   0, 186,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  13,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  64,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 233,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 214,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 115,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 160,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  90,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  92,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  28,   0,   0,   0,   0,   0,   0,   0,   0,   0,  53,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  38,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 128,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 110,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_9  : scenario_type_9 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  31,  31,  31,  30,  31,  29,  31,  28,  31,  27,  31,  26,  31,  25,  31,  24,  31,  23,  31,  22,  31,  21,  31,  20,  31,  19,  31,  18,  31,  17,  31,  16,  31,  15,  31,  14,  31,  13,  31,  12,  31,  11,  31,  10,  31,   9,  31,   8,  31,   7,  31,   6,  31,   5,  31,   4,  31,   3,  31,   2,  31,   1,  31,   0,  31,   0,  31,   0,  31,   0,  31,   0,  31,   0,  31,   0,  31,   0,  31,   0,  31,   0,  31,   0,  31,   0, 230,  31, 230,  30, 230,  29, 230,  28, 230,  27, 230,  26, 230,  25, 230,  24, 230,  23, 230,  22, 230,  21, 230,  20, 230,  19, 230,  18, 230,  17, 230,  16, 230,  15, 230,  14, 230,  13, 230,  12, 230,  11, 230,  10, 230,   9, 230,   8, 230,   7, 230,   6, 230,   5, 230,   4, 230,   3, 230,   2, 230,   1, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0,  33,  31,  33,  30,  33,  29,  33,  28,  33,  27,  33,  26,  33,  25,  33,  24,  33,  23,  33,  22,  33,  21,  33,  20,  33,  19,  33,  18,  33,  17,  33,  16,  33,  15,  33,  14,  33,  13,  33,  12,  33,  11,  33,  10,  33,   9,  33,   8,  33,   7,  33,   6,  33,   5,  33,   4,  33,   3,  33,   2,  33,   1,  33,   0,  33,   0,  33,   0,  33,   0,  33,   0,  33,   0,  33,   0,  33,   0,  33,   0,  33,   0,  33,   0,  33,   0,  33,   0,  33,   0,  33,   0,  33,   0,  33,   0,  21,  31,  21,  30,  21,  29,  21,  28,  21,  27,  21,  26,  21,  25,  21,  24,  21,  23,  21,  22,  21,  21,  21,  20,  21,  19,  21,  18,  21,  17,  21,  16,  21,  15,  21,  14,  21,  13,  21,  12,  21,  11,  21,  10,  21,   9,  21,   8,  21,   7,  21,   6,  87,  31,  87,  30,  87,  29,  87,  28,  87,  27,  87,  26,  87,  25,  87,  24,  87,  23,  87,  22,  87,  21,  87,  20,  87,  19,  87,  18,  87,  17, 200,  31, 200,  30, 200,  29, 200,  28, 200,  27, 200,  26, 200,  25, 200,  24, 200,  23, 200,  22, 200,  21, 200,  20, 200,  19, 200,  18, 200,  17, 200,  16, 200,  15, 200,  14, 200,  13, 200,  12, 200,  11, 200,  10, 200,   9, 200,   8, 200,   7, 200,   6, 200,   5, 200,   4, 200,   3, 200,   2, 200,   1, 200,   0,  58,  31,  58,  30,  58,  29,  58,  28,  58,  27,  58,  26,  58,  25,  58,  24,  58,  23,  58,  22,  58,  21,  58,  20,  58,  19,  58,  18,  58,  17,  58,  16,  58,  15,  58,  14,  58,  13,  58,  12,  58,  11,  58,  10,  58,   9,  58,   8,  58,   7,  58,   6,  58,   5,  58,   4,  58,   3,  58,   2, 152,  31, 152,  30, 152,  29, 152,  28, 152,  27, 152,  26, 129,  31, 129,  30, 129,  29, 129,  28, 129,  27, 129,  26, 129,  25, 228,  31, 228,  30, 228,  29, 228,  28, 228,  27, 228,  26, 228,  25, 228,  24, 228,  23, 228,  22, 228,  21, 228,  20, 228,  19, 228,  18, 228,  17, 228,  16, 228,  15, 228,  14, 228,  13, 228,  12, 228,  11, 228,  10, 228,   9, 228,   8, 228,   7, 228,   6, 228,   5, 228,   4, 228,   3, 228,   2, 228,   1, 228,   0, 228,   0, 228,   0, 228,   0, 228,   0, 228,   0, 228,   0, 228,   0, 228,   0, 228,   0, 228,   0, 228,   0, 228,   0, 228,   0, 228,   0, 228,   0, 228,   0, 228,   0, 228,   0, 228,   0, 228,   0, 228,   0, 228,   0,   6,  31,   6,  30,   6,  29,   6,  28,   6,  27,   6,  26,   6,  25,   6,  24,   6,  23,   6,  22,   6,  21,   6,  20,   6,  19,   6,  18,   6,  17,   6,  16,   6,  15,   6,  14,   6,  13,   6,  12,   6,  11,   6,  10,   6,   9,   6,   8,   6,   7,   6,   6,   6,   5,   6,   4,   6,   3,   6,   2,   6,   1,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0, 250,  31, 250,  30, 250,  29, 250,  28, 250,  27, 250,  26, 250,  25, 250,  24, 250,  23, 250,  22, 250,  21, 250,  20, 250,  19, 250,  18, 250,  17, 250,  16, 250,  15, 250,  14, 250,  13, 250,  12, 250,  11, 250,  10, 250,   9, 250,   8, 250,   7, 250,   6, 250,   5, 250,   4, 250,   3, 250,   2, 250,   1, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 179,  31, 179,  30, 179,  29, 179,  28, 179,  27, 179,  26, 179,  25, 179,  24, 179,  23, 179,  22, 179,  21, 179,  20, 179,  19, 179,  18, 179,  17, 179,  16, 179,  15, 179,  14, 179,  13, 179,  12, 179,  11, 179,  10, 179,   9, 179,   8, 179,   7, 179,   6, 179,   5, 179,   4, 179,   3, 179,   2, 179,   1, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 151,  31, 151,  30, 151,  29, 151,  28, 151,  27, 151,  26, 151,  25, 151,  24, 151,  23, 151,  22, 151,  21, 151,  20, 151,  19, 151,  18, 151,  17, 151,  16, 241,  31, 241,  30, 241,  29, 241,  28, 241,  27, 241,  26, 241,  25, 241,  24, 241,  23, 241,  22, 241,  21, 241,  20, 241,  19, 241,  18, 241,  17, 241,  16, 241,  15, 241,  14, 241,  13, 241,  12, 241,  11, 241,  10, 241,   9, 241,   8, 241,   7, 241,   6, 241,   5, 241,   4, 241,   3, 241,   2, 241,   1, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 133,  31, 133,  30, 186,  31, 186,  30, 186,  29, 186,  28, 186,  27, 186,  26, 186,  25, 186,  24, 186,  23, 186,  22, 186,  21, 186,  20, 186,  19, 186,  18, 186,  17, 186,  16, 186,  15,  13,  31,  13,  30,  13,  29,  13,  28,  13,  27,  13,  26,  13,  25,  64,  31,  64,  30,  64,  29,  64,  28,  64,  27,  64,  26,  64,  25,  64,  24,  64,  23,  64,  22,  64,  21,  64,  20,  64,  19,  64,  18,  64,  17,  64,  16,  64,  15,  64,  14,  64,  13,  64,  12,  64,  11,  64,  10,  64,   9,  64,   8,  64,   7,  64,   6,  64,   5,  64,   4,  64,   3,  64,   2,  64,   1,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0, 233,  31, 233,  30, 233,  29, 233,  28, 233,  27, 233,  26, 233,  25, 233,  24, 233,  23, 233,  22, 233,  21, 233,  20, 214,  31, 214,  30, 214,  29, 214,  28, 214,  27, 214,  26, 214,  25, 214,  24, 214,  23, 214,  22, 214,  21, 214,  20, 214,  19, 214,  18, 214,  17, 214,  16, 214,  15, 214,  14, 214,  13, 214,  12, 214,  11, 214,  10, 214,   9, 214,   8, 214,   7, 214,   6, 214,   5, 214,   4, 214,   3, 115,  31, 115,  30, 115,  29, 115,  28, 115,  27, 115,  26, 115,  25, 115,  24, 115,  23, 115,  22, 115,  21, 115,  20, 115,  19, 115,  18, 115,  17, 115,  16, 115,  15, 115,  14, 115,  13, 115,  12, 115,  11, 115,  10, 115,   9, 115,   8, 115,   7, 115,   6, 115,   5, 115,   4, 115,   3, 115,   2, 115,   1, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 160,  31, 160,  30, 160,  29, 160,  28, 160,  27, 160,  26,  90,  31,  90,  30,  90,  29,  90,  28,  90,  27,  90,  26,  90,  25,  90,  24,  90,  23,  90,  22,  90,  21,  90,  20,  90,  19,  90,  18,  90,  17,  90,  16,  90,  15,  90,  14,  90,  13,  90,  12,  90,  11,  90,  10,  90,   9,  90,   8,  90,   7,  90,   6,  90,   5,  90,   4,  90,   3,  90,   2,  90,   1,  90,   0,  90,   0,  90,   0,  90,   0,  90,   0,  90,   0,  90,   0,  90,   0,  90,   0,  90,   0,  90,   0,  90,   0,  90,   0,  90,   0,  90,   0,  90,   0,  90,   0,  90,   0,  90,   0,  90,   0,  90,   0,  90,   0,  92,  31,  92,  30,  92,  29,  92,  28,  92,  27,  92,  26,  92,  25,  92,  24,  92,  23,  92,  22,  92,  21,  92,  20,  92,  19,  92,  18,  92,  17,  92,  16,  92,  15,  92,  14,  92,  13,  92,  12,  92,  11,  92,  10,  92,   9,  92,   8,  92,   7,  92,   6,  92,   5,  92,   4,  92,   3,  92,   2,  92,   1,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  92,   0,  28,  31,  28,  30,  28,  29,  28,  28,  28,  27,  53,  31,  53,  30,  53,  29,  53,  28,  53,  27,  53,  26,  53,  25,  53,  24,  53,  23,  53,  22,  53,  21,  53,  20,  53,  19,  53,  18,  53,  17,  53,  16,  53,  15,  53,  14,  53,  13,  53,  12,  53,  11,  53,  10,  53,   9,  53,   8,  53,   7,  53,   6,  53,   5,  53,   4,  53,   3,  53,   2,  38,  31,  38,  30,  38,  29,  38,  28,  38,  27,  38,  26,  38,  25,  38,  24,  38,  23,  38,  22,  38,  21,  38,  20,  38,  19,  38,  18,  38,  17,  38,  16,  38,  15,  38,  14,  38,  13,  38,  12,  38,  11,  38,  10,  38,   9,  38,   8,  38,   7,  38,   6,  38,   5,  38,   4,  38,   3,  38,   2,  38,   1, 128,  31, 128,  30, 128,  29, 128,  28, 128,  27, 128,  26, 128,  25, 128,  24, 128,  23, 128,  22, 128,  21, 128,  20, 128,  19, 128,  18, 128,  17, 128,  16, 128,  15, 128,  14, 128,  13, 128,  12, 128,  11, 128,  10, 128,   9, 128,   8, 128,   7, 128,   6, 128,   5, 110,  31, 110,  30, 110,  29, 110,  28, 110,  27, 110,  26, 110,  25, 110,  24, 110,  23, 110,  22, 110,  21, 110,  20, 110,  19, 110,  18, 110,  17, 110,  16, 110,  15, 110,  14, 110,  13);
	constant SCENARIO_ADDRESS_9 : integer := 18437;


	--Scenario 10
	constant SCENARIO_LENGTH_10 : integer := 1022;
	type scenario_type_10 is array (0 to SCENARIO_LENGTH_10*2-1) of integer;
	signal scenario_input_10 : scenario_type_10 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 120,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 109,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  16,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  51,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 173,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 119,   0,   0,   0,   0,   0, 122,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   6,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 120,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   7,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 224,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 243,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  86,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  35,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  60,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 104,   0,   0,   0,   0,   0, 170,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  52,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 134,   0,   0,   0,   0,   0, 185,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 222,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 231,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_10  : scenario_type_10 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 120,  31, 120,  30, 120,  29, 120,  28, 120,  27, 120,  26, 120,  25, 120,  24, 120,  23, 120,  22, 120,  21, 120,  20, 120,  19, 120,  18, 120,  17, 120,  16, 120,  15, 120,  14, 120,  13, 120,  12, 120,  11, 120,  10, 120,   9, 120,   8, 120,   7, 120,   6, 120,   5, 120,   4, 120,   3, 120,   2, 120,   1, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 109,  31, 109,  30, 109,  29, 109,  28, 109,  27, 109,  26, 109,  25, 109,  24, 109,  23, 109,  22, 109,  21, 109,  20, 109,  19, 109,  18, 109,  17, 109,  16,  16,  31,  16,  30,  16,  29,  16,  28,  16,  27,  16,  26,  16,  25,  16,  24,  16,  23,  16,  22,  16,  21,  16,  20,  16,  19,  16,  18,  16,  17,  16,  16,  16,  15,  16,  14,  16,  13,  16,  12,  16,  11,  16,  10,  16,   9,  16,   8,  16,   7,  16,   6,  16,   5,  16,   4,  16,   3,  16,   2,  16,   1,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  51,  31,  51,  30,  51,  29,  51,  28,  51,  27,  51,  26,  51,  25,  51,  24,  51,  23,  51,  22,  51,  21,  51,  20,  51,  19,  51,  18,  51,  17,  51,  16,  51,  15,  51,  14,  51,  13,  51,  12,  51,  11,  51,  10,  51,   9,  51,   8, 173,  31, 173,  30, 173,  29, 173,  28, 173,  27, 173,  26, 173,  25, 173,  24, 173,  23, 173,  22, 173,  21, 173,  20, 173,  19, 173,  18, 173,  17, 173,  16, 173,  15, 173,  14, 119,  31, 119,  30, 119,  29, 122,  31, 122,  30, 122,  29, 122,  28, 122,  27, 122,  26, 122,  25, 122,  24, 122,  23, 122,  22, 122,  21, 122,  20, 122,  19, 122,  18, 122,  17, 122,  16, 122,  15, 122,  14, 122,  13, 122,  12, 122,  11, 122,  10, 122,   9, 122,   8, 122,   7, 122,   6, 122,   5, 122,   4, 122,   3, 122,   2, 122,   1, 122,   0, 122,   0, 122,   0,   6,  31,   6,  30,   6,  29,   6,  28,   6,  27,   6,  26,   6,  25,   6,  24,   6,  23,   6,  22,   6,  21,   6,  20,   6,  19,   6,  18,   6,  17,   6,  16,   6,  15,   6,  14,   6,  13,   6,  12,   6,  11,   6,  10,   6,   9,   6,   8,   6,   7,   6,   6,   6,   5,   6,   4,   6,   3,   6,   2,   6,   1,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0, 120,  31, 120,  30, 120,  29, 120,  28, 120,  27, 120,  26, 120,  25, 120,  24, 120,  23, 120,  22, 120,  21, 120,  20, 120,  19, 120,  18, 120,  17, 120,  16, 120,  15, 120,  14, 120,  13, 120,  12, 120,  11, 120,  10, 120,   9, 120,   8, 120,   7, 120,   6, 120,   5, 120,   4, 120,   3, 120,   2, 120,   1, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0,   7,  31,   7,  30,   7,  29,   7,  28,   7,  27,   7,  26,   7,  25,   7,  24,   7,  23,   7,  22,   7,  21,   7,  20,   7,  19,   7,  18,   7,  17,   7,  16,   7,  15,   7,  14,   7,  13,   7,  12,   7,  11,   7,  10,   7,   9,   7,   8,   7,   7,   7,   6,   7,   5,   7,   4,   7,   3,   7,   2,   7,   1,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0, 224,  31, 224,  30, 224,  29, 224,  28, 224,  27, 224,  26, 224,  25, 224,  24, 224,  23, 224,  22, 224,  21, 224,  20, 224,  19, 224,  18, 224,  17, 224,  16, 224,  15, 224,  14, 224,  13, 224,  12, 224,  11, 224,  10, 224,   9, 224,   8, 224,   7, 224,   6, 224,   5, 224,   4, 224,   3, 224,   2, 224,   1, 224,   0, 224,   0, 224,   0, 243,  31, 243,  30, 243,  29, 243,  28, 243,  27, 243,  26, 243,  25, 243,  24, 243,  23, 243,  22, 243,  21, 243,  20, 243,  19, 243,  18,  86,  31,  86,  30,  86,  29,  86,  28,  86,  27,  86,  26,  86,  25,  86,  24,  86,  23,  86,  22,  86,  21,  86,  20,  86,  19,  86,  18,  86,  17,  86,  16,  86,  15,  86,  14,  86,  13,  86,  12,  86,  11,  35,  31,  35,  30,  35,  29,  35,  28,  35,  27,  35,  26,  35,  25,  35,  24,  35,  23,  35,  22,  35,  21,  35,  20,  35,  19,  35,  18,  35,  17,  35,  16,  35,  15,  35,  14,  35,  13,  35,  12,  35,  11,  35,  10,  35,   9,  35,   8,  35,   7,  35,   6,  35,   5,  35,   4,  35,   3,  35,   2,  60,  31,  60,  30,  60,  29,  60,  28,  60,  27,  60,  26,  60,  25,  60,  24,  60,  23,  60,  22,  60,  21,  60,  20,  60,  19,  60,  18,  60,  17,  60,  16,  60,  15,  60,  14,  60,  13,  60,  12,  60,  11,  60,  10,  60,   9,  60,   8,  60,   7,  60,   6,  60,   5,  60,   4,  60,   3,  60,   2,  60,   1,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0, 104,  31, 104,  30, 104,  29, 170,  31, 170,  30, 170,  29, 170,  28, 170,  27, 170,  26, 170,  25, 170,  24, 170,  23, 170,  22, 170,  21, 170,  20, 170,  19, 170,  18, 170,  17, 170,  16, 170,  15, 170,  14, 170,  13, 170,  12, 170,  11, 170,  10, 170,   9, 170,   8, 170,   7, 170,   6, 170,   5, 170,   4, 170,   3, 170,   2, 170,   1, 170,   0, 170,   0, 170,   0, 170,   0, 170,   0, 170,   0, 170,   0,  52,  31,  52,  30,  52,  29,  52,  28,  52,  27,  52,  26,  52,  25,  52,  24,  52,  23,  52,  22,  52,  21,  52,  20,  52,  19,  52,  18,  52,  17,  52,  16,  52,  15,  52,  14,  52,  13,  52,  12,  52,  11,  52,  10,  52,   9,  52,   8,  52,   7,  52,   6,  52,   5,  52,   4,  52,   3,  52,   2,  52,   1,  52,   0,  52,   0,  52,   0,  52,   0,  52,   0,  52,   0,  52,   0,  52,   0,  52,   0,  52,   0,  52,   0,  52,   0,  52,   0, 134,  31, 134,  30, 134,  29, 185,  31, 185,  30, 185,  29, 185,  28, 185,  27, 185,  26, 185,  25, 185,  24, 185,  23, 185,  22, 185,  21, 185,  20, 185,  19, 185,  18, 185,  17, 185,  16, 185,  15, 185,  14, 185,  13, 185,  12, 185,  11, 185,  10, 185,   9, 185,   8, 185,   7, 185,   6, 185,   5, 185,   4, 185,   3, 185,   2, 185,   1, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 222,  31, 222,  30, 222,  29, 222,  28, 222,  27, 222,  26, 222,  25, 222,  24, 222,  23, 222,  22, 222,  21, 222,  20, 222,  19, 222,  18, 222,  17, 222,  16, 222,  15, 222,  14, 222,  13, 222,  12, 222,  11, 231,  31, 231,  30, 231,  29, 231,  28, 231,  27, 231,  26, 231,  25, 231,  24, 231,  23, 231,  22, 231,  21, 231,  20, 231,  19, 231,  18, 231,  17, 231,  16, 231,  15, 231,  14, 231,  13, 231,  12, 231,  11, 231,  10, 231,   9, 231,   8, 231,   7, 231,   6, 231,   5, 231,   4, 231,   3, 231,   2, 231,   1, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0, 231,   0);
	constant SCENARIO_ADDRESS_10 : integer := 20484;


	--Scenario 11
	constant SCENARIO_LENGTH_11 : integer := 988;
	type scenario_type_11 is array (0 to SCENARIO_LENGTH_11*2-1) of integer;
	signal scenario_input_11 : scenario_type_11 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 196,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  78,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  17,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 210,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 247,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  96,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  41,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 245,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  89,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 228,   0,   0,   0,  69,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 239,   0,   0,   0, 189,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 246,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 198,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 102,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 175,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  83,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  18,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 194,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 228,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 149,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 104,   0,   0,   0,   0,   0,   0,   0,   0,   0, 110,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 218,   0, 156,   0,  36,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 160,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 246,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 209,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_11  : scenario_type_11 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 196,  31, 196,  30, 196,  29, 196,  28, 196,  27, 196,  26, 196,  25, 196,  24, 196,  23, 196,  22, 196,  21, 196,  20, 196,  19, 196,  18, 196,  17, 196,  16, 196,  15, 196,  14, 196,  13, 196,  12, 196,  11, 196,  10, 196,   9, 196,   8, 196,   7, 196,   6, 196,   5, 196,   4, 196,   3, 196,   2, 196,   1, 196,   0, 196,   0, 196,   0, 196,   0, 196,   0, 196,   0, 196,   0, 196,   0, 196,   0, 196,   0, 196,   0, 196,   0, 196,   0, 196,   0, 196,   0, 196,   0,  78,  31,  78,  30,  78,  29,  78,  28,  78,  27,  78,  26,  78,  25,  78,  24,  78,  23,  78,  22,  78,  21,  78,  20,  78,  19,  78,  18,  78,  17,  78,  16,  78,  15,  78,  14,  78,  13,  78,  12,  78,  11,  78,  10,  78,   9,  78,   8,  78,   7,  78,   6,  78,   5,  78,   4,  78,   3,  78,   2,  78,   1,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  17,  31,  17,  30,  17,  29,  17,  28,  17,  27,  17,  26,  17,  25,  17,  24,  17,  23,  17,  22,  17,  21,  17,  20,  17,  19,  17,  18,  17,  17,  17,  16,  17,  15,  17,  14,  17,  13,  17,  12,  17,  11,  17,  10,  17,   9,  17,   8,  17,   7,  17,   6,  17,   5,  17,   4,  17,   3,  17,   2,  17,   1,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0, 210,  31, 210,  30, 210,  29, 210,  28, 210,  27, 210,  26, 210,  25, 210,  24, 210,  23, 210,  22, 247,  31, 247,  30, 247,  29, 247,  28, 247,  27, 247,  26, 247,  25, 247,  24, 247,  23, 247,  22,  96,  31,  96,  30,  96,  29,  96,  28,  96,  27,  96,  26,  96,  25,  96,  24,  96,  23,  96,  22,  96,  21,  96,  20,  96,  19,  96,  18,  96,  17,  96,  16,  96,  15,  96,  14,  96,  13,  96,  12,  96,  11,  96,  10,  96,   9,  96,   8,  96,   7,  96,   6,  96,   5,  96,   4,  96,   3,  96,   2,  96,   1,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  96,   0,  41,  31,  41,  30,  41,  29,  41,  28,  41,  27,  41,  26,  41,  25,  41,  24,  41,  23,  41,  22,  41,  21,  41,  20,  41,  19,  41,  18,  41,  17,  41,  16,  41,  15,  41,  14,  41,  13,  41,  12,  41,  11,  41,  10,  41,   9,  41,   8,  41,   7,  41,   6,  41,   5,  41,   4,  41,   3,  41,   2,  41,   1,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0,  41,   0, 245,  31, 245,  30, 245,  29, 245,  28, 245,  27, 245,  26, 245,  25, 245,  24, 245,  23,  89,  31,  89,  30,  89,  29,  89,  28,  89,  27,  89,  26,  89,  25,  89,  24,  89,  23,  89,  22,  89,  21,  89,  20,  89,  19,  89,  18,  89,  17,  89,  16,  89,  15,  89,  14,  89,  13,  89,  12,  89,  11,  89,  10,  89,   9,  89,   8,  89,   7,  89,   6,  89,   5,  89,   4,  89,   3,  89,   2,  89,   1,  89,   0,  89,   0,  89,   0,  89,   0,  89,   0,  89,   0,  89,   0,  89,   0,  89,   0,  89,   0,  89,   0,  89,   0, 228,  31, 228,  30,  69,  31,  69,  30,  69,  29,  69,  28,  69,  27,  69,  26,  69,  25,  69,  24, 239,  31, 239,  30, 189,  31, 189,  30, 189,  29, 189,  28, 189,  27, 189,  26, 189,  25, 189,  24, 189,  23, 189,  22, 189,  21, 189,  20, 189,  19, 189,  18, 189,  17, 189,  16, 189,  15, 189,  14, 189,  13, 189,  12, 189,  11, 189,  10, 189,   9, 189,   8, 189,   7, 189,   6, 189,   5, 189,   4, 189,   3, 189,   2, 189,   1, 189,   0, 189,   0, 246,  31, 246,  30, 246,  29, 246,  28, 246,  27, 246,  26, 246,  25, 246,  24, 246,  23, 246,  22, 246,  21, 246,  20, 246,  19, 246,  18, 246,  17, 246,  16, 246,  15, 246,  14, 246,  13, 246,  12, 246,  11, 246,  10, 246,   9, 246,   8, 246,   7, 246,   6, 246,   5, 246,   4, 246,   3, 246,   2, 246,   1, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 246,   0, 198,  31, 198,  30, 198,  29, 198,  28, 198,  27, 198,  26, 198,  25, 198,  24, 198,  23, 198,  22, 198,  21, 198,  20, 198,  19, 198,  18, 198,  17, 198,  16, 198,  15, 198,  14, 198,  13, 198,  12, 198,  11, 198,  10, 198,   9, 198,   8, 198,   7, 198,   6, 102,  31, 102,  30, 102,  29, 102,  28, 102,  27, 102,  26, 102,  25, 102,  24, 102,  23, 102,  22, 102,  21, 102,  20, 102,  19, 102,  18, 102,  17, 102,  16, 102,  15, 102,  14, 175,  31, 175,  30, 175,  29, 175,  28, 175,  27, 175,  26, 175,  25, 175,  24, 175,  23, 175,  22, 175,  21, 175,  20, 175,  19, 175,  18, 175,  17, 175,  16, 175,  15, 175,  14, 175,  13, 175,  12, 175,  11, 175,  10, 175,   9, 175,   8, 175,   7, 175,   6, 175,   5, 175,   4, 175,   3, 175,   2, 175,   1, 175,   0, 175,   0, 175,   0, 175,   0,  83,  31,  83,  30,  83,  29,  83,  28,  83,  27,  83,  26,  83,  25,  83,  24,  83,  23,  83,  22,  83,  21,  83,  20,  83,  19,  83,  18,  83,  17,  83,  16,  83,  15,  83,  14,  83,  13,  83,  12,  83,  11,  83,  10,  83,   9,  83,   8,  83,   7,  83,   6,  83,   5,  83,   4,  83,   3,  83,   2,  83,   1,  83,   0,  83,   0,  83,   0,  83,   0,  18,  31,  18,  30,  18,  29,  18,  28,  18,  27,  18,  26,  18,  25,  18,  24,  18,  23,  18,  22,  18,  21,  18,  20,  18,  19,  18,  18,  18,  17,  18,  16,  18,  15,  18,  14,  18,  13,  18,  12, 194,  31, 194,  30, 194,  29, 194,  28, 194,  27, 194,  26, 228,  31, 228,  30, 228,  29, 228,  28, 228,  27, 228,  26, 228,  25, 228,  24, 228,  23, 228,  22, 228,  21, 228,  20, 228,  19, 228,  18, 228,  17, 228,  16, 228,  15, 228,  14, 228,  13, 228,  12, 228,  11, 228,  10, 149,  31, 149,  30, 149,  29, 149,  28, 149,  27, 149,  26, 149,  25, 149,  24, 149,  23, 149,  22, 149,  21, 149,  20, 149,  19, 149,  18, 149,  17, 149,  16, 149,  15, 149,  14, 149,  13, 149,  12, 149,  11, 149,  10, 149,   9, 149,   8, 149,   7, 149,   6, 149,   5, 149,   4, 149,   3, 149,   2, 149,   1, 104,  31, 104,  30, 104,  29, 104,  28, 104,  27, 110,  31, 110,  30, 110,  29, 110,  28, 110,  27, 110,  26, 218,  31, 156,  31,  36,  31,  36,  30,  36,  29,  36,  28,  36,  27,  36,  26,  36,  25,  36,  24,  36,  23,  36,  22,  36,  21,  36,  20,  36,  19,  36,  18,  36,  17,  36,  16,  36,  15,  36,  14,  36,  13,  36,  12,  36,  11,  36,  10,  36,   9,  36,   8,  36,   7,  36,   6,  36,   5,  36,   4,  36,   3,  36,   2,  36,   1,  36,   0,  36,   0,  36,   0,  36,   0,  36,   0,  36,   0,  36,   0,  36,   0,  36,   0,  36,   0,  36,   0,  36,   0, 160,  31, 160,  30, 160,  29, 160,  28, 160,  27, 160,  26, 160,  25, 160,  24, 160,  23, 160,  22, 160,  21, 160,  20, 160,  19, 160,  18, 160,  17, 160,  16, 160,  15, 246,  31, 246,  30, 246,  29, 246,  28, 246,  27, 246,  26, 246,  25, 246,  24, 246,  23, 246,  22, 246,  21, 246,  20, 246,  19, 246,  18, 246,  17, 246,  16, 246,  15, 246,  14, 209,  31, 209,  30, 209,  29, 209,  28, 209,  27);
	constant SCENARIO_ADDRESS_11 : integer := 22558;


	--Scenario 12
	constant SCENARIO_LENGTH_12 : integer := 1015;
	type scenario_type_12 is array (0 to SCENARIO_LENGTH_12*2-1) of integer;
	signal scenario_input_12 : scenario_type_12 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 209,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 135,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 144,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 227,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 105,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 230,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 237,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  19,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 214,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 205,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  68,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 166,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 177,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 194,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 150,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  62,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 135,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 123,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 173,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 194,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   3,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 255,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 101,   0,   0,   0,  82,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 207,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 120,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  67,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  21,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  21,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_12  : scenario_type_12 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 209,  31, 209,  30, 209,  29, 209,  28, 209,  27, 209,  26, 209,  25, 209,  24, 209,  23, 209,  22, 209,  21, 209,  20, 209,  19, 209,  18, 209,  17, 209,  16, 209,  15, 209,  14, 209,  13, 209,  12, 209,  11, 209,  10, 209,   9, 209,   8, 209,   7, 209,   6, 209,   5, 209,   4, 209,   3, 209,   2, 209,   1, 209,   0, 209,   0, 209,   0, 209,   0, 209,   0, 209,   0, 209,   0, 209,   0, 209,   0, 209,   0, 209,   0, 209,   0, 135,  31, 135,  30, 135,  29, 135,  28, 135,  27, 135,  26, 135,  25, 135,  24, 135,  23, 135,  22, 135,  21, 135,  20, 135,  19, 135,  18, 135,  17, 135,  16, 135,  15, 135,  14, 135,  13, 135,  12, 135,  11, 135,  10, 135,   9, 135,   8, 135,   7, 135,   6, 135,   5, 135,   4, 135,   3, 135,   2, 144,  31, 144,  30, 144,  29, 144,  28, 144,  27, 144,  26, 144,  25, 144,  24, 144,  23, 144,  22, 144,  21, 144,  20, 144,  19, 144,  18, 144,  17, 144,  16, 227,  31, 227,  30, 227,  29, 227,  28, 227,  27, 227,  26, 227,  25, 227,  24, 227,  23, 227,  22, 227,  21, 227,  20, 227,  19, 227,  18, 227,  17, 227,  16, 227,  15, 227,  14, 227,  13, 105,  31, 105,  30, 105,  29, 105,  28, 105,  27, 105,  26, 105,  25, 230,  31, 230,  30, 230,  29, 230,  28, 230,  27, 230,  26, 230,  25, 230,  24, 230,  23, 230,  22, 230,  21, 230,  20, 230,  19, 230,  18, 230,  17, 230,  16, 230,  15, 230,  14, 230,  13, 230,  12, 230,  11, 230,  10, 230,   9, 230,   8, 230,   7, 230,   6, 230,   5, 230,   4, 230,   3, 230,   2, 230,   1, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 230,   0, 237,  31, 237,  30, 237,  29, 237,  28, 237,  27, 237,  26, 237,  25, 237,  24, 237,  23, 237,  22, 237,  21, 237,  20, 237,  19, 237,  18, 237,  17, 237,  16, 237,  15, 237,  14, 237,  13, 237,  12, 237,  11, 237,  10, 237,   9, 237,   8, 237,   7, 237,   6, 237,   5, 237,   4, 237,   3, 237,   2, 237,   1, 237,   0, 237,   0, 237,   0, 237,   0, 237,   0, 237,   0, 237,   0, 237,   0, 237,   0, 237,   0, 237,   0,  19,  31,  19,  30,  19,  29,  19,  28,  19,  27,  19,  26,  19,  25,  19,  24,  19,  23,  19,  22,  19,  21,  19,  20,  19,  19,  19,  18,  19,  17,  19,  16,  19,  15,  19,  14,  19,  13,  19,  12,  19,  11,  19,  10,  19,   9,  19,   8,  19,   7,  19,   6,  19,   5,  19,   4,  19,   3,  19,   2,  19,   1,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0, 214,  31, 214,  30, 214,  29, 214,  28, 214,  27, 214,  26, 214,  25, 214,  24, 214,  23, 214,  22, 205,  31, 205,  30, 205,  29, 205,  28, 205,  27, 205,  26, 205,  25, 205,  24, 205,  23, 205,  22, 205,  21, 205,  20, 205,  19, 205,  18, 205,  17, 205,  16, 205,  15, 205,  14, 205,  13, 205,  12, 205,  11, 205,  10, 205,   9, 205,   8, 205,   7, 205,   6, 205,   5, 205,   4, 205,   3, 205,   2, 205,   1, 205,   0, 205,   0, 205,   0, 205,   0, 205,   0,  68,  31,  68,  30,  68,  29,  68,  28,  68,  27,  68,  26,  68,  25,  68,  24,  68,  23,  68,  22,  68,  21,  68,  20,  68,  19,  68,  18,  68,  17,  68,  16,  68,  15,  68,  14,  68,  13,  68,  12,  68,  11,  68,  10,  68,   9,  68,   8,  68,   7,  68,   6,  68,   5,  68,   4,  68,   3,  68,   2,  68,   1,  68,   0,  68,   0,  68,   0,  68,   0,  68,   0,  68,   0,  68,   0,  68,   0,  68,   0,  68,   0,  68,   0,  68,   0,  68,   0,  68,   0,  68,   0,  68,   0,  68,   0,  68,   0,  68,   0,  68,   0, 166,  31, 166,  30, 166,  29, 166,  28, 166,  27, 166,  26, 166,  25, 166,  24, 166,  23, 166,  22, 166,  21, 166,  20, 166,  19, 166,  18, 166,  17, 166,  16, 166,  15, 166,  14, 166,  13, 166,  12, 166,  11, 166,  10, 166,   9, 166,   8, 166,   7, 166,   6, 166,   5, 166,   4, 166,   3, 166,   2, 166,   1, 177,  31, 177,  30, 177,  29, 177,  28, 177,  27, 177,  26, 177,  25, 177,  24, 177,  23, 177,  22, 177,  21, 177,  20, 177,  19, 177,  18, 177,  17, 177,  16, 177,  15, 177,  14, 177,  13, 177,  12, 177,  11, 177,  10, 177,   9, 177,   8, 177,   7, 194,  31, 194,  30, 194,  29, 194,  28, 194,  27, 194,  26, 194,  25, 194,  24, 194,  23, 194,  22, 194,  21, 194,  20, 194,  19, 194,  18, 194,  17, 194,  16, 194,  15, 194,  14, 194,  13, 194,  12, 194,  11, 194,  10, 194,   9, 194,   8, 194,   7, 194,   6, 194,   5, 194,   4, 194,   3, 194,   2, 194,   1, 150,  31, 150,  30, 150,  29, 150,  28, 150,  27, 150,  26, 150,  25, 150,  24, 150,  23, 150,  22, 150,  21, 150,  20, 150,  19, 150,  18, 150,  17, 150,  16, 150,  15, 150,  14, 150,  13, 150,  12, 150,  11, 150,  10, 150,   9, 150,   8, 150,   7, 150,   6, 150,   5, 150,   4, 150,   3, 150,   2, 150,   1, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0,  62,  31,  62,  30,  62,  29,  62,  28,  62,  27,  62,  26,  62,  25,  62,  24,  62,  23,  62,  22,  62,  21,  62,  20,  62,  19,  62,  18,  62,  17,  62,  16,  62,  15,  62,  14,  62,  13,  62,  12,  62,  11,  62,  10,  62,   9,  62,   8,  62,   7,  62,   6,  62,   5,  62,   4,  62,   3,  62,   2,  62,   1,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0,  62,   0, 135,  31, 135,  30, 135,  29, 135,  28, 135,  27, 135,  26, 135,  25, 135,  24, 135,  23, 135,  22, 135,  21, 135,  20, 135,  19, 135,  18, 135,  17, 135,  16, 135,  15, 123,  31, 123,  30, 123,  29, 123,  28, 123,  27, 123,  26, 123,  25, 123,  24, 123,  23, 123,  22, 123,  21, 123,  20, 123,  19, 123,  18, 123,  17, 173,  31, 173,  30, 173,  29, 173,  28, 173,  27, 173,  26, 194,  31, 194,  30, 194,  29, 194,  28, 194,  27, 194,  26, 194,  25, 194,  24,   3,  31,   3,  30,   3,  29,   3,  28,   3,  27,   3,  26,   3,  25,   3,  24,   3,  23, 255,  31, 255,  30, 255,  29, 255,  28, 255,  27, 255,  26, 255,  25, 255,  24, 255,  23, 255,  22, 255,  21, 255,  20, 255,  19, 255,  18, 255,  17, 255,  16, 255,  15, 255,  14, 255,  13, 255,  12, 255,  11, 255,  10, 255,   9, 255,   8, 255,   7, 255,   6, 255,   5, 255,   4, 255,   3, 255,   2, 255,   1, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 101,  31, 101,  30,  82,  31,  82,  30,  82,  29,  82,  28,  82,  27,  82,  26,  82,  25,  82,  24,  82,  23,  82,  22,  82,  21,  82,  20,  82,  19,  82,  18,  82,  17,  82,  16,  82,  15,  82,  14,  82,  13,  82,  12,  82,  11,  82,  10,  82,   9,  82,   8,  82,   7,  82,   6,  82,   5,  82,   4,  82,   3,  82,   2,  82,   1,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0,  82,   0, 207,  31, 207,  30, 207,  29, 207,  28, 207,  27, 207,  26, 207,  25, 207,  24, 207,  23, 207,  22, 207,  21, 207,  20, 207,  19, 207,  18, 207,  17, 207,  16, 207,  15, 207,  14, 207,  13, 207,  12, 207,  11, 207,  10, 207,   9, 207,   8, 207,   7, 207,   6, 207,   5, 207,   4, 207,   3, 207,   2, 207,   1, 207,   0, 207,   0, 207,   0, 207,   0, 207,   0, 207,   0, 207,   0, 207,   0, 207,   0, 207,   0, 207,   0, 207,   0, 207,   0, 207,   0, 207,   0, 207,   0, 207,   0, 207,   0, 207,   0, 207,   0, 207,   0, 207,   0, 207,   0, 207,   0, 120,  31, 120,  30, 120,  29, 120,  28, 120,  27, 120,  26, 120,  25, 120,  24, 120,  23, 120,  22, 120,  21, 120,  20, 120,  19, 120,  18, 120,  17, 120,  16, 120,  15, 120,  14, 120,  13, 120,  12,  67,  31,  67,  30,  67,  29,  67,  28,  67,  27,  67,  26,  67,  25,  67,  24,  67,  23,  67,  22,  67,  21,  67,  20,  67,  19,  67,  18,  67,  17,  67,  16,  67,  15,  67,  14,  67,  13,  67,  12,  67,  11,  67,  10,  67,   9,  67,   8,  67,   7,  67,   6,  67,   5,  67,   4,  67,   3,  67,   2,  67,   1,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  21,  31,  21,  30,  21,  29,  21,  28,  21,  27,  21,  26,  21,  25,  21,  24,  21,  23,  21,  22,  21,  21,  21,  20,  21,  19,  21,  18,  21,  17,  21,  16,  21,  15,  21,  14,  21,  13,  21,  12,  21,  11,  21,  10,  21,   9,  21,   8,  21,   7,  21,   6,  21,   5,  21,   4,  21,   3,  21,   2,  21,   1,  21,  31,  21,  30,  21,  29,  21,  28,  21,  27,  21,  26,  21,  25,  21,  24,  21,  23,  21,  22,  21,  21);
	constant SCENARIO_ADDRESS_12 : integer := 24583;


	--Scenario 13
	constant SCENARIO_LENGTH_13 : integer := 1001;
	type scenario_type_13 is array (0 to SCENARIO_LENGTH_13*2-1) of integer;
	signal scenario_input_13 : scenario_type_13 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  60,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  24,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  11,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 197,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  91,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  74,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  99,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 132,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 206,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  32,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 205,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 142,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   2,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 113,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 119,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 173,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 219,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  58,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 119,   0,   0,   0, 239,   0,   0,   0,   0,   0,   0,   0, 146,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 234,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  85,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  96,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 189,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   6,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_13  : scenario_type_13 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  60,  31,  60,  30,  60,  29,  60,  28,  60,  27,  60,  26,  60,  25,  60,  24,  60,  23,  60,  22,  60,  21,  60,  20,  60,  19,  60,  18,  60,  17,  60,  16,  60,  15,  60,  14,  60,  13,  60,  12,  60,  11,  60,  10,  60,   9,  60,   8,  60,   7,  60,   6,  60,   5,  60,   4,  60,   3,  60,   2,  60,   1,  60,   0,  24,  31,  24,  30,  24,  29,  24,  28,  24,  27,  24,  26,  24,  25,  24,  24,  24,  23,  24,  22,  24,  21,  24,  20,  24,  19,  24,  18,  24,  17,  24,  16,  24,  15,  24,  14,  24,  13,  24,  12,  24,  11,  11,  31,  11,  30,  11,  29,  11,  28,  11,  27,  11,  26,  11,  25,  11,  24,  11,  23,  11,  22,  11,  21,  11,  20,  11,  19,  11,  18,  11,  17,  11,  16,  11,  15,  11,  14,  11,  13,  11,  12,  11,  11,  11,  10,  11,   9,  11,   8,  11,   7,  11,   6,  11,   5,  11,   4,  11,   3,  11,   2,  11,   1,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0,  11,   0, 197,  31, 197,  30, 197,  29, 197,  28, 197,  27, 197,  26, 197,  25, 197,  24, 197,  23, 197,  22, 197,  21, 197,  20, 197,  19, 197,  18, 197,  17, 197,  16, 197,  15, 197,  14, 197,  13, 197,  12, 197,  11, 197,  10, 197,   9, 197,   8, 197,   7, 197,   6, 197,   5, 197,   4, 197,   3, 197,   2, 197,   1, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0,  91,  31,  91,  30,  91,  29,  91,  28,  91,  27,  91,  26,  91,  25,  91,  24,  91,  23,  91,  22,  91,  21,  91,  20,  91,  19,  91,  18,  91,  17,  91,  16,  91,  15,  91,  14,  91,  13,  91,  12,  91,  11,  91,  10,  91,   9,  91,   8,  91,   7,  91,   6,  91,   5,  91,   4,  91,   3,  91,   2,  91,   1,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  74,  31,  74,  30,  74,  29,  74,  28,  74,  27,  74,  26,  74,  25,  74,  24,  74,  23,  74,  22,  74,  21,  74,  20,  74,  19,  99,  31,  99,  30,  99,  29,  99,  28,  99,  27,  99,  26,  99,  25,  99,  24,  99,  23,  99,  22,  99,  21,  99,  20,  99,  19,  99,  18,  99,  17,  99,  16,  99,  15,  99,  14,  99,  13,  99,  12,  99,  11,  99,  10,  99,   9,  99,   8,  99,   7,  99,   6,  99,   5,  99,   4,  99,   3,  99,   2,  99,   1,  99,   0,  99,   0, 132,  31, 132,  30, 132,  29, 132,  28, 132,  27, 132,  26, 132,  25, 132,  24, 132,  23, 132,  22, 132,  21, 132,  20, 132,  19, 132,  18, 132,  17, 132,  16, 132,  15, 132,  14, 132,  13, 132,  12, 206,  31, 206,  30, 206,  29, 206,  28, 206,  27, 206,  26,  32,  31,  32,  30,  32,  29,  32,  28,  32,  27,  32,  26,  32,  25,  32,  24,  32,  23,  32,  22,  32,  21,  32,  20,  32,  19,  32,  18,  32,  17, 205,  31, 205,  30, 205,  29, 205,  28, 205,  27, 205,  26, 205,  25, 205,  24, 205,  23, 205,  22, 205,  21, 205,  20, 205,  19, 205,  18, 205,  17, 205,  16, 205,  15, 205,  14, 205,  13, 205,  12, 205,  11, 205,  10, 205,   9, 205,   8, 205,   7, 205,   6, 205,   5, 205,   4, 205,   3, 205,   2, 205,   1, 205,   0, 205,   0, 205,   0, 205,   0, 205,   0, 205,   0, 205,   0, 142,  31, 142,  30, 142,  29, 142,  28, 142,  27, 142,  26, 142,  25, 142,  24, 142,  23, 142,  22, 142,  21, 142,  20, 142,  19, 142,  18, 142,  17, 142,  16, 142,  15, 142,  14, 142,  13, 142,  12, 142,  11, 142,  10, 142,   9, 142,   8, 142,   7, 142,   6, 142,   5, 142,   4, 142,   3, 142,   2, 142,   1, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0,   2,  31,   2,  30,   2,  29,   2,  28,   2,  27,   2,  26,   2,  25,   2,  24,   2,  23,   2,  22,   2,  21,   2,  20,   2,  19,   2,  18,   2,  17,   2,  16,   2,  15,   2,  14,   2,  13,   2,  12,   2,  11,   2,  10,   2,   9,   2,   8,   2,   7,   2,   6,   2,   5,   2,   4,   2,   3,   2,   2,   2,   1,   2,   0,   2,   0,   2,   0,   2,   0,   2,   0,   2,   0, 113,  31, 113,  30, 113,  29, 113,  28, 113,  27, 113,  26, 113,  25, 113,  24, 113,  23, 113,  22, 113,  21, 113,  20, 113,  19, 113,  18, 113,  17, 113,  16, 113,  15, 113,  14, 113,  13, 113,  12, 113,  11, 113,  10, 113,   9, 113,   8, 113,   7, 113,   6, 113,   5, 113,   4, 113,   3, 113,   2, 113,   1, 113,   0, 113,   0, 113,   0, 113,   0, 113,   0, 113,   0, 113,   0, 113,   0, 113,   0, 119,  31, 119,  30, 119,  29, 119,  28, 119,  27, 119,  26, 119,  25, 119,  24, 119,  23, 119,  22, 119,  21, 119,  20, 119,  19, 173,  31, 173,  30, 173,  29, 173,  28, 173,  27, 173,  26, 173,  25, 173,  24, 173,  23, 173,  22, 173,  21, 173,  20, 173,  19, 173,  18, 173,  17, 173,  16, 173,  15, 173,  14, 173,  13, 173,  12, 173,  11, 173,  10, 173,   9, 173,   8, 173,   7, 173,   6, 173,   5, 173,   4, 173,   3, 173,   2, 173,   1, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 219,  31, 219,  30, 219,  29, 219,  28, 219,  27, 219,  26, 219,  25, 219,  24, 219,  23, 219,  22, 219,  21, 219,  20, 219,  19, 219,  18, 219,  17, 219,  16, 219,  15, 219,  14,  58,  31,  58,  30,  58,  29,  58,  28,  58,  27,  58,  26,  58,  25,  58,  24,  58,  23,  58,  22,  58,  21,  58,  20,  58,  19,  58,  18,  58,  17,  58,  16,  58,  15,  58,  14,  58,  13,  58,  12,  58,  11,  58,  10,  58,   9,  58,   8,  58,   7,  58,   6,  58,   5,  58,   4,  58,   3,  58,   2,  58,   1,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0, 119,  31, 119,  30, 239,  31, 239,  30, 239,  29, 239,  28, 146,  31, 146,  30, 146,  29, 146,  28, 146,  27, 146,  26, 146,  25, 146,  24, 146,  23, 146,  22, 146,  21, 146,  20, 146,  19, 146,  18, 146,  17, 146,  16, 146,  15, 146,  14, 146,  13, 146,  12, 146,  11, 146,  10, 146,   9, 146,   8, 146,   7, 146,   6, 146,   5, 146,   4, 146,   3, 146,   2, 146,   1, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 234,  31, 234,  30, 234,  29, 234,  28, 234,  27, 234,  26, 234,  25, 234,  24, 234,  23, 234,  22, 234,  21, 234,  20, 234,  19, 234,  18, 234,  17, 234,  16, 234,  15, 234,  14, 234,  13, 234,  12, 234,  11, 234,  10, 234,   9, 234,   8, 234,   7, 234,   6, 234,   5, 234,   4, 234,   3, 234,   2, 234,   1, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0, 234,   0,  85,  31,  85,  30,  85,  29,  85,  28,  85,  27,  85,  26,  85,  25,  85,  24,  85,  23,  85,  22,  85,  21,  85,  20,  85,  19,  85,  18,  85,  17,  85,  16,  85,  15,  85,  14,  85,  13,  85,  12,  85,  11,  85,  10,  85,   9,  85,   8,  85,   7,  85,   6,  85,   5,  85,   4,  85,   3,  85,   2,  85,   1,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  85,   0,  96,  31,  96,  30,  96,  29,  96,  28,  96,  27,  96,  26,  96,  25,  96,  24,  96,  23,  96,  22,  96,  21,  96,  20,  96,  19,  96,  18,  96,  17,  96,  16,  96,  15, 189,  31, 189,  30, 189,  29, 189,  28, 189,  27, 189,  26, 189,  25, 189,  24, 189,  23, 189,  22,   6,  31,   6,  30,   6,  29,   6,  28,   6,  27,   6,  26,   6,  25,   6,  24,   6,  23,   6,  22,   6,  21,   6,  20,   6,  19,   6,  18,   6,  17,   6,  16,   6,  15,   6,  14,   6,  13,   6,  12,   6,  11,   6,  10,   6,   9,   6,   8,   6,   7,   6,   6,   6,   5,   6,   4,   6,   3,   6,   2,   6,   1,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0);
	constant SCENARIO_ADDRESS_13 : integer := 26669;


	--Scenario 14
	constant SCENARIO_LENGTH_14 : integer := 1016;
	type scenario_type_14 is array (0 to SCENARIO_LENGTH_14*2-1) of integer;
	signal scenario_input_14 : scenario_type_14 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  99,   0,   0,   0,   0,   0,   0,   0,   0,   0,  34,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  94,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  51,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 222,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   4,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 180,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 204,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 130,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 237,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  20,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 161,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 172,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  11,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  99,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 250,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 135,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  51,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  16,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 144,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 173,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  97,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 205,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 255,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 244,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_14  : scenario_type_14 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  99,  31,  99,  30,  99,  29,  99,  28,  99,  27,  34,  31,  34,  30,  34,  29,  34,  28,  34,  27,  34,  26,  34,  25,  34,  24,  34,  23,  34,  22,  34,  21,  34,  20,  34,  19,  34,  18,  34,  17,  34,  16,  34,  15,  34,  14,  34,  13,  34,  12,  34,  11,  34,  10,  34,   9,  34,   8,  34,   7,  34,   6,  34,   5,  34,   4,  34,   3,  94,  31,  94,  30,  94,  29,  94,  28,  94,  27,  94,  26,  94,  25,  94,  24,  94,  23,  94,  22,  94,  21,  94,  20,  94,  19,  94,  18,  94,  17,  94,  16,  94,  15,  94,  14,  94,  13,  94,  12,  94,  11,  94,  10,  94,   9,  94,   8,  94,   7,  94,   6,  94,   5,  94,   4,  94,   3,  51,  31,  51,  30,  51,  29,  51,  28,  51,  27,  51,  26,  51,  25,  51,  24,  51,  23,  51,  22,  51,  21,  51,  20,  51,  19,  51,  18,  51,  17,  51,  16,  51,  15,  51,  14,  51,  13,  51,  12,  51,  11,  51,  10,  51,   9,  51,   8,  51,   7,  51,   6,  51,   5,  51,   4,  51,   3,  51,   2,  51,   1,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0, 222,  31, 222,  30, 222,  29, 222,  28, 222,  27, 222,  26, 222,  25, 222,  24, 222,  23, 222,  22, 222,  21, 222,  20, 222,  19, 222,  18, 222,  17, 222,  16, 222,  15, 222,  14, 222,  13, 222,  12, 222,  11, 222,  10, 222,   9, 222,   8, 222,   7, 222,   6, 222,   5, 222,   4, 222,   3, 222,   2, 222,   1, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0,   4,  31,   4,  30,   4,  29,   4,  28,   4,  27,   4,  26,   4,  25,   4,  24,   4,  23,   4,  22,   4,  21,   4,  20,   4,  19,   4,  18,   4,  17,   4,  16,   4,  15,   4,  14,   4,  13,   4,  12,   4,  11,   4,  10,   4,   9,   4,   8,   4,   7,   4,   6,   4,   5,   4,   4,   4,   3,   4,   2,   4,   1,   4,   0,   4,   0,   4,   0,   4,   0,   4,   0,   4,   0,   4,   0,   4,   0,   4,   0,   4,   0, 180,  31, 180,  30, 180,  29, 180,  28, 180,  27, 180,  26, 180,  25, 180,  24, 180,  23, 180,  22, 180,  21, 180,  20, 180,  19, 180,  18, 180,  17, 180,  16, 180,  15, 180,  14, 180,  13, 180,  12, 180,  11, 180,  10, 180,   9, 180,   8, 180,   7, 180,   6, 180,   5, 180,   4, 180,   3, 180,   2, 180,   1, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 204,  31, 204,  30, 204,  29, 204,  28, 204,  27, 204,  26, 204,  25, 204,  24, 204,  23, 204,  22, 204,  21, 204,  20, 204,  19, 204,  18, 204,  17, 204,  16, 204,  15, 204,  14, 204,  13, 204,  12, 204,  11, 204,  10, 204,   9, 204,   8, 204,   7, 204,   6, 204,   5, 204,   4, 204,   3, 204,   2, 204,   1, 204,   0, 130,  31, 130,  30, 130,  29, 130,  28, 130,  27, 130,  26, 130,  25, 130,  24, 130,  23, 130,  22, 130,  21, 130,  20, 130,  19, 130,  18, 130,  17, 130,  16, 130,  15, 130,  14, 130,  13, 130,  12, 130,  11, 130,  10, 130,   9, 130,   8, 130,   7, 130,   6, 130,   5, 130,   4, 130,   3, 130,   2, 130,   1, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 237,  31, 237,  30, 237,  29, 237,  28, 237,  27, 237,  26, 237,  25, 237,  24, 237,  23, 237,  22, 237,  21, 237,  20, 237,  19, 237,  18, 237,  17, 237,  16, 237,  15, 237,  14, 237,  13, 237,  12, 237,  11, 237,  10, 237,   9, 237,   8, 237,   7, 237,   6, 237,   5, 237,   4, 237,   3,  20,  31,  20,  30,  20,  29,  20,  28,  20,  27,  20,  26,  20,  25,  20,  24,  20,  23,  20,  22,  20,  21,  20,  20,  20,  19,  20,  18,  20,  17, 161,  31, 161,  30, 161,  29, 161,  28, 161,  27, 161,  26, 161,  25, 161,  24, 161,  23, 161,  22, 161,  21, 161,  20, 161,  19, 161,  18, 161,  17, 161,  16, 161,  15, 161,  14, 161,  13, 161,  12, 161,  11, 161,  10, 161,   9, 161,   8, 161,   7, 161,   6, 161,   5, 161,   4, 161,   3, 161,   2, 161,   1, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 161,   0, 172,  31, 172,  30, 172,  29, 172,  28, 172,  27, 172,  26, 172,  25, 172,  24, 172,  23, 172,  22, 172,  21, 172,  20, 172,  19, 172,  18, 172,  17, 172,  16, 172,  15, 172,  14, 172,  13, 172,  12, 172,  11, 172,  10, 172,   9, 172,   8, 172,   7, 172,   6, 172,   5, 172,   4, 172,   3, 172,   2, 172,   1, 172,   0, 172,   0, 172,   0, 172,   0, 172,   0, 172,   0, 172,   0, 172,   0,  11,  31,  11,  30,  11,  29,  11,  28,  11,  27,  11,  26,  11,  25,  11,  24,  11,  23,  11,  22,  11,  21,  11,  20,  11,  19,  11,  18,  11,  17,  11,  16,  11,  15,  11,  14,  11,  13,  11,  12,  11,  11,  11,  10,  11,   9,  99,  31,  99,  30,  99,  29,  99,  28,  99,  27,  99,  26, 250,  31, 250,  30, 250,  29, 250,  28, 250,  27, 250,  26, 250,  25, 250,  24, 250,  23, 250,  22, 250,  21, 250,  20, 250,  19, 250,  18, 135,  31, 135,  30, 135,  29, 135,  28, 135,  27, 135,  26, 135,  25, 135,  24, 135,  23, 135,  22, 135,  21, 135,  20, 135,  19, 135,  18, 135,  17, 135,  16, 135,  15, 135,  14, 135,  13, 135,  12, 135,  11, 135,  10, 135,   9, 135,   8, 135,   7, 135,   6, 135,   5, 135,   4, 135,   3, 135,   2, 135,   1, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0,  51,  31,  51,  30,  51,  29,  51,  28,  51,  27,  51,  26,  51,  25,  51,  24,  51,  23,  51,  22,  51,  21,  51,  20,  51,  19,  51,  18,  51,  17,  51,  16,  51,  15,  51,  14,  51,  13,  51,  12,  51,  11,  51,  10,  51,   9,  51,   8,  51,   7,  51,   6,  51,   5,  51,   4,  51,   3,  51,   2,  51,   1,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  16,  31,  16,  30,  16,  29,  16,  28,  16,  27,  16,  26,  16,  25,  16,  24,  16,  23,  16,  22,  16,  21,  16,  20,  16,  19,  16,  18,  16,  17,  16,  16,  16,  15,  16,  14,  16,  13,  16,  12,  16,  11,  16,  10,  16,   9,  16,   8,  16,   7,  16,   6,  16,   5,  16,   4,  16,   3,  16,   2,  16,   1,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0, 144,  31, 144,  30, 144,  29, 144,  28, 144,  27, 144,  26, 144,  25, 144,  24, 144,  23, 144,  22, 144,  21, 144,  20, 144,  19, 144,  18, 144,  17, 144,  16, 144,  15, 144,  14, 144,  13, 144,  12, 144,  11, 144,  10, 144,   9, 144,   8, 144,   7, 144,   6, 144,   5, 144,   4, 144,   3, 144,   2, 144,   1, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 144,   0, 173,  31, 173,  30, 173,  29, 173,  28, 173,  27, 173,  26, 173,  25, 173,  24, 173,  23, 173,  22, 173,  21, 173,  20, 173,  19, 173,  18, 173,  17, 173,  16, 173,  15, 173,  14, 173,  13, 173,  12, 173,  11, 173,  10, 173,   9, 173,   8, 173,   7, 173,   6, 173,   5, 173,   4, 173,   3, 173,   2, 173,   1, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0,  97,  31,  97,  30,  97,  29,  97,  28,  97,  27,  97,  26,  97,  25,  97,  24,  97,  23,  97,  22,  97,  21,  97,  20,  97,  19,  97,  18,  97,  17,  97,  16,  97,  15,  97,  14,  97,  13,  97,  12,  97,  11,  97,  10,  97,   9,  97,   8,  97,   7,  97,   6,  97,   5,  97,   4,  97,   3,  97,   2,  97,   1,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0,  97,   0, 205,  31, 205,  30, 205,  29, 205,  28, 205,  27, 205,  26, 205,  25, 205,  24, 205,  23, 205,  22, 205,  21, 205,  20, 205,  19, 205,  18, 255,  31, 255,  30, 255,  29, 255,  28, 255,  27, 255,  26, 255,  25, 255,  24, 255,  23, 255,  22, 255,  21, 255,  20, 255,  19, 255,  18, 255,  17, 255,  16, 255,  15, 255,  14, 255,  13, 255,  12, 255,  11, 255,  10, 255,   9, 255,   8, 255,   7, 255,   6, 255,   5, 255,   4, 255,   3, 255,   2, 255,   1, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 255,   0, 244,  31, 244,  30, 244,  29, 244,  28, 244,  27, 244,  26, 244,  25, 244,  24, 244,  23, 244,  22, 244,  21, 244,  20, 244,  19, 244,  18, 244,  17, 244,  16, 244,  15, 244,  14, 244,  13, 244,  12, 244,  11, 244,  10, 244,   9, 244,   8, 244,   7, 244,   6, 244,   5, 244,   4, 244,   3, 244,   2, 244,   1, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0);
	constant SCENARIO_ADDRESS_14 : integer := 28681;


	--Scenario 15
	constant SCENARIO_LENGTH_15 : integer := 988;
	type scenario_type_15 is array (0 to SCENARIO_LENGTH_15*2-1) of integer;
	signal scenario_input_15 : scenario_type_15 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  93,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 146,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 131,   0, 180,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 165,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 179,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 176,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 139,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  84,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 197,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 214,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 142,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 195,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 186,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 217,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 146,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 141,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 177,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 219,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  16,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 220,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_15  : scenario_type_15 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  93,  31,  93,  30,  93,  29,  93,  28,  93,  27,  93,  26,  93,  25,  93,  24,  93,  23,  93,  22,  93,  21,  93,  20,  93,  19,  93,  18,  93,  17,  93,  16,  93,  15,  93,  14,  93,  13,  93,  12,  93,  11,  93,  10,  93,   9,  93,   8,  93,   7,  93,   6,  93,   5,  93,   4,  93,   3,  93,   2,  93,   1,  93,   0,  93,   0,  93,   0,  93,   0,  93,   0,  93,   0,  93,   0,  93,   0,  93,   0,  93,   0,  93,   0,  93,   0,  93,   0,  93,   0,  93,   0,  93,   0,  93,   0,  93,   0, 146,  31, 146,  30, 146,  29, 146,  28, 146,  27, 146,  26, 146,  25, 146,  24, 146,  23, 146,  22, 146,  21, 146,  20, 146,  19, 146,  18, 146,  17, 146,  16, 146,  15, 146,  14, 146,  13, 146,  12, 146,  11, 146,  10, 146,   9, 146,   8, 131,  31, 180,  31, 180,  30, 180,  29, 180,  28, 180,  27, 180,  26, 180,  25, 180,  24, 180,  23, 180,  22, 180,  21, 180,  20, 180,  19, 180,  18, 180,  17, 180,  16, 180,  15, 180,  14, 180,  13, 165,  31, 165,  30, 165,  29, 165,  28, 165,  27, 165,  26, 165,  25, 165,  24, 165,  23, 165,  22, 165,  21, 165,  20, 165,  19, 165,  18, 165,  17, 165,  16, 165,  15, 165,  14, 165,  13, 165,  12, 165,  11, 165,  10, 165,   9, 165,   8, 165,   7, 165,   6, 165,   5, 165,   4, 165,   3, 165,   2, 165,   1, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 179,  31, 179,  30, 179,  29, 179,  28, 179,  27, 179,  26, 179,  25, 179,  24, 179,  23, 179,  22, 179,  21, 179,  20, 179,  19, 179,  18, 179,  17, 179,  16, 179,  15, 179,  14, 179,  13, 179,  12, 179,  11, 179,  10, 179,   9, 179,   8, 179,   7, 179,   6, 179,   5, 179,   4, 179,   3, 179,   2, 179,   1, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 176,  31, 176,  30, 176,  29, 176,  28, 176,  27, 176,  26, 176,  25, 176,  24, 176,  23, 176,  22, 176,  21, 176,  20, 176,  19, 139,  31, 139,  30, 139,  29, 139,  28, 139,  27, 139,  26, 139,  25, 139,  24, 139,  23, 139,  22, 139,  21, 139,  20, 139,  19, 139,  18, 139,  17, 139,  16, 139,  15, 139,  14, 139,  13, 139,  12, 139,  11, 139,  10, 139,   9, 139,   8, 139,   7, 139,   6, 139,   5, 139,   4, 139,   3, 139,   2, 139,   1, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0,  84,  31,  84,  30,  84,  29,  84,  28,  84,  27,  84,  26,  84,  25,  84,  24,  84,  23,  84,  22,  84,  21,  84,  20,  84,  19,  84,  18,  84,  17,  84,  16,  84,  15,  84,  14,  84,  13,  84,  12,  84,  11,  84,  10,  84,   9,  84,   8, 197,  31, 197,  30, 197,  29, 197,  28, 197,  27, 197,  26, 197,  25, 197,  24, 197,  23, 197,  22, 197,  21, 197,  20, 197,  19, 197,  18, 197,  17, 197,  16, 197,  15, 197,  14, 197,  13, 197,  12, 197,  11, 197,  10, 197,   9, 197,   8, 197,   7, 197,   6, 197,   5, 197,   4, 197,   3, 197,   2, 197,   1, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 214,  31, 214,  30, 214,  29, 214,  28, 214,  27, 214,  26, 214,  25, 214,  24, 214,  23, 214,  22, 214,  21, 214,  20, 214,  19, 214,  18, 214,  17, 214,  16, 214,  15, 214,  14, 214,  13, 214,  12, 214,  11, 214,  10, 214,   9, 214,   8, 214,   7, 214,   6, 214,   5, 214,   4, 214,   3, 214,   2, 214,   1, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 142,  31, 142,  30, 142,  29, 142,  28, 142,  27, 142,  26, 142,  25, 142,  24, 142,  23, 142,  22, 142,  21, 142,  20, 142,  19, 142,  18, 142,  17, 142,  16, 142,  15, 142,  14, 142,  13, 142,  12, 142,  11, 142,  10, 142,   9, 142,   8, 142,   7, 142,   6, 142,   5, 142,   4, 142,   3, 142,   2, 142,   1, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 195,  31, 195,  30, 195,  29, 195,  28, 195,  27, 195,  26, 195,  25, 195,  24, 195,  23, 195,  22, 195,  21, 195,  20, 195,  19, 195,  18, 195,  17, 195,  16, 195,  15, 195,  14, 195,  13, 195,  12, 195,  11, 195,  10, 195,   9, 195,   8, 195,   7, 195,   6, 195,   5, 195,   4, 195,   3, 195,   2, 195,   1, 195,   0, 195,   0, 195,   0, 195,   0, 195,   0, 195,   0, 195,   0, 195,   0, 195,   0, 195,   0, 186,  31, 186,  30, 186,  29, 186,  28, 186,  27, 186,  26, 186,  25, 186,  24, 186,  23, 186,  22, 186,  21, 186,  20, 186,  19, 186,  18, 186,  17, 186,  16, 186,  15, 186,  14, 186,  13, 186,  12, 186,  11, 186,  10, 186,   9, 186,   8, 186,   7, 186,   6, 186,   5, 186,   4, 186,   3, 186,   2, 186,   1, 186,   0, 186,   0, 186,   0, 186,   0, 186,   0, 217,  31, 217,  30, 217,  29, 217,  28, 217,  27, 217,  26, 217,  25, 217,  24, 217,  23, 217,  22, 217,  21, 217,  20, 217,  19, 217,  18, 217,  17, 217,  16, 217,  15, 217,  14, 217,  13, 217,  12, 217,  11, 217,  10, 217,   9, 217,   8, 217,   7, 217,   6, 217,   5, 217,   4, 217,   3, 217,   2, 217,   1, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 217,   0, 146,  31, 146,  30, 146,  29, 146,  28, 146,  27, 146,  26, 146,  25, 146,  24, 146,  23, 146,  22, 146,  21, 146,  20, 146,  19, 146,  18, 146,  17, 146,  16, 146,  15, 146,  14, 146,  13, 146,  12, 141,  31, 141,  30, 141,  29, 141,  28, 141,  27, 141,  26, 141,  25, 141,  24, 141,  23, 141,  22, 141,  21, 141,  20, 141,  19, 141,  18, 141,  17, 141,  16, 141,  15, 141,  14, 141,  13, 141,  12, 141,  11, 141,  10, 141,   9, 141,   8, 141,   7, 141,   6, 141,   5, 141,   4, 141,   3, 141,   2, 141,   1, 141,   0, 141,   0, 141,   0, 141,   0, 141,   0, 141,   0, 141,   0, 141,   0, 141,   0, 177,  31, 177,  30, 177,  29, 177,  28, 177,  27, 177,  26, 177,  25, 219,  31, 219,  30, 219,  29, 219,  28, 219,  27, 219,  26, 219,  25, 219,  24, 219,  23, 219,  22, 219,  21, 219,  20, 219,  19, 219,  18, 219,  17, 219,  16, 219,  15, 219,  14, 219,  13, 219,  12,  16,  31,  16,  30,  16,  29,  16,  28,  16,  27,  16,  26,  16,  25,  16,  24,  16,  23,  16,  22,  16,  21,  16,  20,  16,  19,  16,  18,  16,  17,  16,  16,  16,  15,  16,  14,  16,  13,  16,  12, 220,  31, 220,  30, 220,  29, 220,  28, 220,  27, 220,  26, 220,  25, 220,  24, 220,  23, 220,  22, 220,  21, 220,  20, 220,  19, 220,  18, 220,  17, 220,  16, 220,  15, 220,  14, 220,  13, 220,  12, 220,  11, 220,  10, 220,   9, 220,   8, 220,   7, 220,   6, 220,   5, 220,   4, 220,   3, 220,   2, 220,   1, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0);
	constant SCENARIO_ADDRESS_15 : integer := 30762;


	--Scenario 16
	constant SCENARIO_LENGTH_16 : integer := 1;
	type scenario_type_16 is array (0 to SCENARIO_LENGTH_16*2-1) of integer;
	signal scenario_input_16 : scenario_type_16 := (7,   7);
	signal scenario_full_16  : scenario_type_16 := (7,   7);
	constant SCENARIO_ADDRESS_16 : integer := 33519;
	--This sequence is going to be ignored by the component
	--as the i_k parameter is will be set to zero


	--Scenario 17
	constant SCENARIO_LENGTH_17 : integer := 1011;
	type scenario_type_17 is array (0 to SCENARIO_LENGTH_17*2-1) of integer;
	signal scenario_input_17 : scenario_type_17 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 217,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 204,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   5,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 162,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 132,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  63,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  27,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 103,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  63,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  58,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 223,   0,   0,   0,   0,   0, 111,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 206,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 103,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 149,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  35,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 168,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 178,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 165,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 251,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   9,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  12,   0,   0,   0,   0,   0,   0,   0, 204,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  16,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_17  : scenario_type_17 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 217,  31, 217,  30, 217,  29, 217,  28, 217,  27, 217,  26, 217,  25, 217,  24, 217,  23, 217,  22, 217,  21, 217,  20, 217,  19, 217,  18, 217,  17, 217,  16, 217,  15, 217,  14, 217,  13, 217,  12, 217,  11, 217,  10, 217,   9, 217,   8, 204,  31, 204,  30, 204,  29, 204,  28, 204,  27, 204,  26, 204,  25, 204,  24, 204,  23, 204,  22, 204,  21, 204,  20, 204,  19, 204,  18, 204,  17, 204,  16,   5,  31,   5,  30,   5,  29,   5,  28,   5,  27,   5,  26,   5,  25,   5,  24,   5,  23,   5,  22,   5,  21,   5,  20,   5,  19,   5,  18,   5,  17,   5,  16,   5,  15,   5,  14,   5,  13,   5,  12,   5,  11,   5,  10,   5,   9,   5,   8,   5,   7,   5,   6,   5,   5,   5,   4,   5,   3,   5,   2,   5,   1,   5,   0,   5,   0,   5,   0,   5,   0,   5,   0,   5,   0,   5,   0,   5,   0,   5,   0,   5,   0,   5,   0,   5,   0,   5,   0,   5,   0,   5,   0,   5,   0,   5,   0,   5,   0,   5,   0,   5,   0,   5,   0,   5,   0,   5,   0, 162,  31, 162,  30, 162,  29, 162,  28, 162,  27, 162,  26, 162,  25, 162,  24, 162,  23, 162,  22, 162,  21, 162,  20, 162,  19, 162,  18, 162,  17, 162,  16, 162,  15, 162,  14, 162,  13, 162,  12, 162,  11, 162,  10, 162,   9, 162,   8, 162,   7, 162,   6, 162,   5, 162,   4, 162,   3, 162,   2, 162,   1, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 132,  31, 132,  30, 132,  29, 132,  28, 132,  27, 132,  26, 132,  25, 132,  24, 132,  23, 132,  22, 132,  21, 132,  20, 132,  19, 132,  18, 132,  17, 132,  16, 132,  15, 132,  14, 132,  13, 132,  12, 132,  11, 132,  10, 132,   9, 132,   8, 132,   7, 132,   6, 132,   5, 132,   4, 132,   3, 132,   2, 132,   1, 132,   0, 132,   0, 132,   0, 132,   0, 132,   0, 132,   0, 132,   0, 132,   0, 132,   0, 132,   0, 132,   0, 132,   0,  63,  31,  63,  30,  63,  29,  63,  28,  63,  27,  63,  26,  63,  25,  63,  24,  63,  23,  63,  22,  63,  21,  63,  20,  63,  19,  63,  18,  63,  17,  63,  16,  63,  15,  63,  14,  63,  13,  63,  12,  63,  11,  63,  10,  63,   9,  63,   8,  63,   7,  63,   6,  63,   5,  63,   4,  63,   3,  63,   2,  63,   1,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  27,  31,  27,  30,  27,  29,  27,  28,  27,  27,  27,  26,  27,  25,  27,  24,  27,  23,  27,  22,  27,  21,  27,  20,  27,  19,  27,  18,  27,  17,  27,  16,  27,  15,  27,  14,  27,  13,  27,  12,  27,  11,  27,  10,  27,   9,  27,   8,  27,   7,  27,   6,  27,   5,  27,   4,  27,   3,  27,   2,  27,   1,  27,   0,  27,   0,  27,   0,  27,   0,  27,   0, 103,  31, 103,  30, 103,  29, 103,  28, 103,  27, 103,  26, 103,  25, 103,  24, 103,  23, 103,  22, 103,  21, 103,  20, 103,  19,  63,  31,  63,  30,  63,  29,  63,  28,  63,  27,  63,  26,  63,  25,  63,  24,  63,  23,  63,  22,  63,  21,  63,  20,  63,  19,  63,  18,  63,  17,  63,  16,  63,  15,  63,  14,  63,  13,  63,  12,  63,  11,  63,  10,  63,   9,  63,   8,  63,   7,  63,   6,  63,   5,  63,   4,  63,   3,  63,   2,  63,   1,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  58,  31,  58,  30,  58,  29,  58,  28,  58,  27,  58,  26,  58,  25,  58,  24,  58,  23,  58,  22,  58,  21,  58,  20,  58,  19,  58,  18,  58,  17,  58,  16,  58,  15,  58,  14,  58,  13,  58,  12,  58,  11,  58,  10,  58,   9,  58,   8,  58,   7,  58,   6,  58,   5,  58,   4,  58,   3,  58,   2,  58,   1, 223,  31, 223,  30, 223,  29, 111,  31, 111,  30, 111,  29, 111,  28, 111,  27, 111,  26, 111,  25, 111,  24, 111,  23, 111,  22, 111,  21, 111,  20, 111,  19, 111,  18, 111,  17, 111,  16, 111,  15, 111,  14, 111,  13, 111,  12, 111,  11, 111,  10, 111,   9, 111,   8, 111,   7, 111,   6, 111,   5, 111,   4, 111,   3, 111,   2, 111,   1, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 206,  31, 206,  30, 206,  29, 206,  28, 206,  27, 206,  26, 206,  25, 206,  24, 206,  23, 206,  22, 206,  21, 206,  20, 206,  19, 206,  18, 206,  17, 206,  16, 206,  15, 206,  14, 206,  13, 206,  12, 206,  11, 206,  10, 206,   9, 206,   8, 206,   7, 206,   6, 206,   5, 206,   4, 206,   3, 206,   2, 206,   1, 206,   0, 206,   0, 206,   0, 206,   0, 103,  31, 103,  30, 103,  29, 103,  28, 103,  27, 103,  26, 103,  25, 103,  24, 103,  23, 103,  22, 103,  21, 103,  20, 103,  19, 103,  18, 103,  17, 103,  16, 103,  15, 103,  14, 103,  13, 103,  12, 103,  11, 103,  10, 103,   9, 103,   8, 103,   7, 103,   6, 103,   5, 103,   4, 103,   3, 103,   2, 103,   1, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 149,  31, 149,  30, 149,  29, 149,  28, 149,  27, 149,  26, 149,  25, 149,  24, 149,  23, 149,  22, 149,  21, 149,  20, 149,  19, 149,  18, 149,  17, 149,  16, 149,  15, 149,  14, 149,  13, 149,  12, 149,  11, 149,  10, 149,   9, 149,   8, 149,   7, 149,   6, 149,   5, 149,   4, 149,   3, 149,   2, 149,   1, 149,   0, 149,   0, 149,   0,  35,  31,  35,  30,  35,  29,  35,  28,  35,  27,  35,  26,  35,  25,  35,  24,  35,  23,  35,  22,  35,  21,  35,  20,  35,  19,  35,  18,  35,  17,  35,  16,  35,  15,  35,  14,  35,  13,  35,  12,  35,  11,  35,  10,  35,   9,  35,   8,  35,   7,  35,   6,  35,   5,  35,   4,  35,   3,  35,   2,  35,   1,  35,   0,  35,   0,  35,   0,  35,   0,  35,   0,  35,   0, 168,  31, 168,  30, 168,  29, 168,  28, 168,  27, 168,  26, 168,  25, 168,  24, 168,  23, 168,  22, 168,  21, 168,  20, 168,  19, 168,  18, 168,  17, 168,  16, 168,  15, 168,  14, 168,  13, 168,  12, 168,  11, 168,  10, 168,   9, 168,   8, 168,   7, 168,   6, 168,   5, 168,   4, 168,   3, 168,   2, 168,   1, 168,   0, 168,   0, 168,   0, 168,   0, 168,   0, 168,   0, 168,   0, 168,   0, 168,   0, 168,   0, 168,   0, 168,   0, 168,   0, 168,   0, 168,   0, 168,   0, 168,   0, 168,   0, 168,   0, 168,   0, 178,  31, 178,  30, 178,  29, 178,  28, 178,  27, 178,  26, 178,  25, 178,  24, 178,  23, 178,  22, 178,  21, 178,  20, 178,  19, 178,  18, 178,  17, 178,  16, 178,  15, 178,  14, 178,  13, 178,  12, 178,  11, 178,  10, 178,   9, 178,   8, 165,  31, 165,  30, 165,  29, 165,  28, 165,  27, 165,  26, 165,  25, 165,  24, 165,  23, 165,  22, 165,  21, 165,  20, 165,  19, 165,  18, 165,  17, 165,  16, 165,  15, 165,  14, 165,  13, 165,  12, 165,  11, 165,  10, 165,   9, 165,   8, 165,   7, 165,   6, 165,   5, 165,   4, 165,   3, 165,   2, 165,   1, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 165,   0, 251,  31, 251,  30, 251,  29, 251,  28, 251,  27, 251,  26, 251,  25, 251,  24, 251,  23, 251,  22, 251,  21, 251,  20,   9,  31,   9,  30,   9,  29,   9,  28,   9,  27,   9,  26,   9,  25,   9,  24,   9,  23,   9,  22,   9,  21,   9,  20,   9,  19,   9,  18,   9,  17,   9,  16,   9,  15,   9,  14,   9,  13,   9,  12,   9,  11,   9,  10,   9,   9,   9,   8,   9,   7,   9,   6,   9,   5,   9,   4,   9,   3,   9,   2,   9,   1,   9,   0,   9,   0,   9,   0,   9,   0,   9,   0,   9,   0,   9,   0,   9,   0,   9,   0,   9,   0,   9,   0,   9,   0,   9,   0,  12,  31,  12,  30,  12,  29,  12,  28, 204,  31, 204,  30, 204,  29, 204,  28, 204,  27, 204,  26, 204,  25, 204,  24, 204,  23, 204,  22, 204,  21, 204,  20, 204,  19, 204,  18, 204,  17, 204,  16, 204,  15, 204,  14, 204,  13, 204,  12, 204,  11, 204,  10, 204,   9, 204,   8, 204,   7, 204,   6, 204,   5, 204,   4, 204,   3, 204,   2, 204,   1, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0, 204,   0,  16,  31,  16,  30,  16,  29,  16,  28,  16,  27,  16,  26,  16,  25,  16,  24,  16,  23,  16,  22,  16,  21,  16,  20,  16,  19,  16,  18);
	constant SCENARIO_ADDRESS_17 : integer := 34823;


	--Scenario 18
	constant SCENARIO_LENGTH_18 : integer := 1003;
	type scenario_type_18 is array (0 to SCENARIO_LENGTH_18*2-1) of integer;
	signal scenario_input_18 : scenario_type_18 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 192,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   7,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  25,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 118,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  63,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  63,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  60,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 162,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 143,   0,   0,   0,   0,   0,   0,   0,   0,   0, 245,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 115,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 127,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  56,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 143,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  74,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  13,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 138,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 140,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 111,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 173,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  74,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 228,   0,   0,   0,   0,   0,   0,   0, 186,   0,   0,   0, 160,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  11,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 189,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  15,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 185,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  42,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_18  : scenario_type_18 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 192,  31, 192,  30, 192,  29, 192,  28, 192,  27, 192,  26, 192,  25, 192,  24, 192,  23, 192,  22, 192,  21, 192,  20, 192,  19, 192,  18, 192,  17, 192,  16, 192,  15, 192,  14, 192,  13, 192,  12,   7,  31,   7,  30,   7,  29,   7,  28,   7,  27,   7,  26,   7,  25,   7,  24,   7,  23,   7,  22,   7,  21,   7,  20,  25,  31,  25,  30,  25,  29,  25,  28,  25,  27,  25,  26,  25,  25,  25,  24,  25,  23,  25,  22,  25,  21,  25,  20,  25,  19,  25,  18,  25,  17,  25,  16,  25,  15,  25,  14,  25,  13,  25,  12,  25,  11,  25,  10,  25,   9,  25,   8,  25,   7,  25,   6,  25,   5,  25,   4,  25,   3,  25,   2,  25,   1,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0, 118,  31, 118,  30, 118,  29, 118,  28, 118,  27, 118,  26, 118,  25, 118,  24, 118,  23, 118,  22, 118,  21, 118,  20, 118,  19, 118,  18, 118,  17, 118,  16, 118,  15, 118,  14, 118,  13, 118,  12, 118,  11, 118,  10, 118,   9, 118,   8, 118,   7, 118,   6, 118,   5, 118,   4, 118,   3, 118,   2, 118,   1, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0,  63,  31,  63,  30,  63,  29,  63,  28,  63,  27,  63,  26,  63,  25,  63,  24,  63,  23,  63,  22,  63,  21,  63,  20,  63,  19,  63,  18,  63,  17,  63,  16,  63,  15,  63,  14,  63,  13,  63,  12,  63,  11,  63,  10,  63,   9,  63,   8,  63,   7,  63,   6,  63,   5,  63,   4,  63,   3,  63,   2,  63,   1,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,   0,  63,  31,  63,  30,  63,  29,  63,  28,  63,  27,  63,  26,  63,  25,  63,  24,  63,  23,  63,  22,  63,  21,  63,  20,  63,  19,  63,  18,  63,  17,  63,  16,  63,  15,  63,  14,  63,  13,  63,  12,  60,  31,  60,  30,  60,  29,  60,  28,  60,  27,  60,  26,  60,  25,  60,  24,  60,  23,  60,  22,  60,  21,  60,  20,  60,  19,  60,  18,  60,  17,  60,  16,  60,  15,  60,  14,  60,  13,  60,  12,  60,  11,  60,  10,  60,   9,  60,   8,  60,   7,  60,   6,  60,   5,  60,   4,  60,   3, 162,  31, 162,  30, 162,  29, 162,  28, 162,  27, 162,  26, 162,  25, 162,  24, 162,  23, 162,  22, 162,  21, 162,  20, 162,  19, 162,  18, 162,  17, 162,  16, 162,  15, 162,  14, 162,  13, 162,  12, 162,  11, 162,  10, 162,   9, 162,   8, 162,   7, 162,   6, 162,   5, 162,   4, 162,   3, 162,   2, 162,   1, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 143,  31, 143,  30, 143,  29, 143,  28, 143,  27, 245,  31, 245,  30, 245,  29, 245,  28, 245,  27, 245,  26, 245,  25, 245,  24, 245,  23, 245,  22, 245,  21, 245,  20, 245,  19, 245,  18, 245,  17, 245,  16, 245,  15, 245,  14, 245,  13, 245,  12, 245,  11, 245,  10, 245,   9, 245,   8, 245,   7, 245,   6, 245,   5, 245,   4, 245,   3, 245,   2, 245,   1, 245,   0, 245,   0, 245,   0, 245,   0, 245,   0, 245,   0, 245,   0, 245,   0, 245,   0, 245,   0, 245,   0, 245,   0, 245,   0, 245,   0, 245,   0, 245,   0, 245,   0, 245,   0, 245,   0, 245,   0, 245,   0, 245,   0, 115,  31, 115,  30, 115,  29, 115,  28, 115,  27, 115,  26, 115,  25, 115,  24, 115,  23, 115,  22, 115,  21, 115,  20, 115,  19, 115,  18, 115,  17, 115,  16, 115,  15, 115,  14, 115,  13, 115,  12, 115,  11, 115,  10, 115,   9, 115,   8, 115,   7, 115,   6, 115,   5, 115,   4, 115,   3, 115,   2, 115,   1, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 115,   0, 127,  31, 127,  30, 127,  29, 127,  28, 127,  27, 127,  26, 127,  25, 127,  24, 127,  23, 127,  22, 127,  21, 127,  20, 127,  19, 127,  18, 127,  17, 127,  16, 127,  15, 127,  14, 127,  13, 127,  12, 127,  11, 127,  10, 127,   9, 127,   8, 127,   7, 127,   6,  56,  31,  56,  30,  56,  29,  56,  28,  56,  27,  56,  26,  56,  25,  56,  24,  56,  23,  56,  22,  56,  21,  56,  20,  56,  19,  56,  18,  56,  17,  56,  16,  56,  15,  56,  14,  56,  13,  56,  12,  56,  11,  56,  10,  56,   9,  56,   8,  56,   7,  56,   6,  56,   5,  56,   4,  56,   3,  56,   2, 143,  31, 143,  30, 143,  29, 143,  28, 143,  27, 143,  26, 143,  25, 143,  24, 143,  23, 143,  22, 143,  21, 143,  20, 143,  19, 143,  18, 143,  17, 143,  16, 143,  15, 143,  14, 143,  13, 143,  12, 143,  11, 143,  10, 143,   9, 143,   8, 143,   7, 143,   6, 143,   5, 143,   4, 143,   3, 143,   2, 143,   1, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0,  74,  31,  74,  30,  74,  29,  74,  28,  74,  27,  74,  26,  74,  25,  74,  24,  74,  23,  74,  22,  74,  21,  74,  20,  74,  19,  74,  18,  74,  17,  74,  16,  74,  15,  74,  14,  74,  13,  74,  12,  74,  11,  74,  10,  74,   9,  74,   8,  74,   7,  74,   6,  13,  31,  13,  30,  13,  29,  13,  28,  13,  27,  13,  26,  13,  25,  13,  24,  13,  23,  13,  22,  13,  21,  13,  20,  13,  19,  13,  18,  13,  17,  13,  16,  13,  15,  13,  14,  13,  13,  13,  12,  13,  11,  13,  10,  13,   9,  13,   8,  13,   7,  13,   6,  13,   5,  13,   4,  13,   3,  13,   2,  13,   1,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0,  13,   0, 138,  31, 138,  30, 138,  29, 138,  28, 138,  27, 138,  26, 138,  25, 138,  24, 138,  23, 138,  22, 138,  21, 138,  20, 138,  19, 138,  18, 138,  17, 138,  16, 138,  15, 138,  14, 138,  13, 138,  12, 138,  11, 138,  10, 138,   9, 138,   8, 138,   7, 138,   6, 138,   5, 138,   4, 138,   3, 138,   2, 138,   1, 138,   0, 138,   0, 138,   0, 138,   0, 138,   0, 138,   0, 138,   0, 138,   0, 138,   0, 138,   0, 138,   0, 138,   0, 138,   0, 138,   0, 138,   0, 138,   0, 138,   0, 140,  31, 140,  30, 140,  29, 140,  28, 140,  27, 140,  26, 140,  25, 140,  24, 140,  23, 140,  22, 140,  21, 140,  20, 140,  19, 140,  18, 140,  17, 140,  16, 140,  15, 140,  14, 140,  13, 140,  12, 140,  11, 140,  10, 140,   9, 140,   8, 140,   7, 140,   6, 140,   5, 140,   4, 140,   3, 140,   2, 140,   1, 140,   0, 140,   0, 140,   0, 140,   0, 140,   0, 111,  31, 111,  30, 111,  29, 111,  28, 111,  27, 111,  26, 111,  25, 111,  24, 111,  23, 111,  22, 111,  21, 111,  20, 111,  19, 111,  18, 111,  17, 111,  16, 111,  15, 111,  14, 111,  13, 111,  12, 111,  11, 111,  10, 111,   9, 111,   8, 111,   7, 111,   6, 111,   5, 111,   4, 111,   3, 111,   2, 111,   1, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 111,   0, 173,  31, 173,  30, 173,  29, 173,  28, 173,  27, 173,  26, 173,  25, 173,  24, 173,  23, 173,  22, 173,  21, 173,  20, 173,  19, 173,  18, 173,  17, 173,  16, 173,  15, 173,  14, 173,  13, 173,  12, 173,  11, 173,  10, 173,   9, 173,   8, 173,   7, 173,   6, 173,   5, 173,   4, 173,   3, 173,   2, 173,   1, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0,  74,  31,  74,  30,  74,  29,  74,  28,  74,  27,  74,  26,  74,  25, 228,  31, 228,  30, 228,  29, 228,  28, 186,  31, 186,  30, 160,  31, 160,  30, 160,  29, 160,  28, 160,  27, 160,  26, 160,  25, 160,  24, 160,  23, 160,  22, 160,  21, 160,  20, 160,  19, 160,  18, 160,  17, 160,  16, 160,  15, 160,  14, 160,  13, 160,  12, 160,  11, 160,  10, 160,   9, 160,   8, 160,   7, 160,   6, 160,   5, 160,   4, 160,   3, 160,   2, 160,   1, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0,  11,  31,  11,  30,  11,  29,  11,  28,  11,  27,  11,  26,  11,  25,  11,  24,  11,  23,  11,  22,  11,  21,  11,  20,  11,  19,  11,  18,  11,  17,  11,  16, 189,  31, 189,  30, 189,  29, 189,  28, 189,  27, 189,  26, 189,  25, 189,  24,  15,  31,  15,  30,  15,  29,  15,  28,  15,  27,  15,  26, 185,  31, 185,  30, 185,  29, 185,  28, 185,  27, 185,  26, 185,  25, 185,  24, 185,  23, 185,  22, 185,  21, 185,  20, 185,  19, 185,  18, 185,  17, 185,  16, 185,  15, 185,  14, 185,  13, 185,  12, 185,  11, 185,  10, 185,   9,  42,  31,  42,  30,  42,  29,  42,  28,  42,  27,  42,  26,  42,  25,  42,  24,  42,  23,  42,  22,  42,  21,  42,  20,  42,  19,  42,  18,  42,  17,  42,  16,  42,  15,  42,  14,  42,  13,  42,  12,  42,  11,  42,  10,  42,   9,  42,   8,  42,   7,  42,   6,  42,   5,  42,   4,  42,   3,  42,   2,  42,   1,  42,   0,  42,   0,  42,   0,  42,   0,  42,   0,  42,   0,  42,   0,  42,   0,  42,   0,  42,   0,  42,   0,  42,   0,  42,   0,  42,   0,  42,   0,  42,   0,  42,   0,  42,   0,  42,   0,  42,   0,  42,   0,  42,   0,  42,   0,  42,   0);
	constant SCENARIO_ADDRESS_18 : integer := 36888;


	--Scenario 19
	constant SCENARIO_LENGTH_19 : integer := 996;
	type scenario_type_19 is array (0 to SCENARIO_LENGTH_19*2-1) of integer;
	signal scenario_input_19 : scenario_type_19 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 139,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 107,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 175,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 173,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 155,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 137,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  77,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   5,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 123,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 129,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 208,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 154,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 250,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 242,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 243,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 175,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 210,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 103,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   5,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_19  : scenario_type_19 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 139,  31, 139,  30, 139,  29, 139,  28, 139,  27, 139,  26, 139,  25, 139,  24, 139,  23, 139,  22, 139,  21, 139,  20, 139,  19, 139,  18, 139,  17, 139,  16, 139,  15, 139,  14, 139,  13, 139,  12, 139,  11, 139,  10, 139,   9, 139,   8, 139,   7, 139,   6, 139,   5, 139,   4, 139,   3, 139,   2, 139,   1, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 107,  31, 107,  30, 107,  29, 107,  28, 107,  27, 107,  26, 107,  25, 107,  24, 107,  23, 107,  22, 107,  21, 107,  20, 107,  19, 107,  18, 107,  17, 107,  16, 107,  15, 107,  14, 107,  13, 107,  12, 107,  11, 107,  10, 107,   9, 107,   8, 107,   7, 107,   6, 107,   5, 107,   4, 107,   3, 107,   2, 107,   1, 107,   0, 107,   0, 175,  31, 175,  30, 175,  29, 175,  28, 175,  27, 175,  26, 175,  25, 175,  24, 175,  23, 175,  22, 175,  21, 175,  20, 175,  19, 175,  18, 175,  17, 175,  16, 175,  15, 175,  14, 175,  13, 175,  12, 175,  11, 175,  10, 175,   9, 175,   8, 175,   7, 175,   6, 173,  31, 173,  30, 173,  29, 173,  28, 173,  27, 173,  26, 173,  25, 173,  24, 173,  23, 173,  22, 173,  21, 173,  20, 173,  19, 173,  18, 173,  17, 173,  16, 173,  15, 173,  14, 173,  13, 173,  12, 173,  11, 173,  10, 173,   9, 173,   8, 173,   7, 173,   6, 173,   5, 173,   4, 173,   3, 173,   2, 173,   1, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 173,   0, 155,  31, 155,  30, 155,  29, 155,  28, 155,  27, 155,  26, 155,  25, 155,  24, 137,  31, 137,  30, 137,  29, 137,  28, 137,  27, 137,  26, 137,  25, 137,  24, 137,  23, 137,  22, 137,  21, 137,  20, 137,  19, 137,  18, 137,  17, 137,  16, 137,  15, 137,  14, 137,  13, 137,  12, 137,  11, 137,  10, 137,   9, 137,   8, 137,   7, 137,   6, 137,   5, 137,   4, 137,   3, 137,   2, 137,   1, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0,  77,  31,  77,  30,  77,  29,  77,  28,  77,  27,  77,  26,  77,  25,  77,  24,  77,  23,  77,  22,  77,  21,  77,  20,  77,  19,  77,  18,  77,  17,  77,  16,  77,  15,  77,  14,  77,  13,  77,  12,  77,  11,  77,  10,  77,   9,  77,   8,  77,   7,  77,   6,  77,   5,  77,   4,   5,  31,   5,  30,   5,  29,   5,  28,   5,  27,   5,  26,   5,  25,   5,  24,   5,  23,   5,  22,   5,  21,   5,  20,   5,  19,   5,  18,   5,  17,   5,  16,   5,  15,   5,  14,   5,  13,   5,  12,   5,  11,   5,  10,   5,   9,   5,   8,   5,   7,   5,   6,   5,   5,   5,   4,   5,   3,   5,   2,   5,   1, 123,  31, 123,  30, 123,  29, 123,  28, 123,  27, 123,  26, 123,  25, 123,  24, 123,  23, 123,  22, 123,  21, 123,  20, 123,  19, 123,  18, 123,  17, 123,  16, 123,  15, 123,  14, 123,  13, 123,  12, 123,  11, 123,  10, 123,   9, 123,   8, 123,   7, 123,   6, 123,   5, 123,   4, 123,   3, 123,   2, 123,   1, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 129,  31, 129,  30, 129,  29, 129,  28, 129,  27, 129,  26, 129,  25, 129,  24, 129,  23, 129,  22, 129,  21, 129,  20, 129,  19, 129,  18, 129,  17, 129,  16, 129,  15, 129,  14, 129,  13, 129,  12, 129,  11, 129,  10, 129,   9, 129,   8, 129,   7, 129,   6, 129,   5, 129,   4, 129,   3, 129,   2, 129,   1, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 208,  31, 208,  30, 208,  29, 208,  28, 208,  27, 208,  26, 208,  25, 208,  24, 208,  23, 208,  22, 208,  21, 208,  20, 208,  19, 208,  18, 208,  17, 208,  16, 208,  15, 208,  14, 208,  13, 208,  12, 208,  11, 208,  10, 208,   9, 208,   8, 208,   7, 208,   6, 208,   5, 208,   4, 208,   3, 208,   2, 208,   1, 208,   0, 208,   0, 208,   0, 208,   0, 208,   0, 208,   0, 208,   0, 208,   0, 208,   0, 208,   0, 208,   0, 208,   0, 208,   0, 208,   0, 208,   0, 208,   0, 208,   0, 208,   0, 208,   0, 208,   0, 154,  31, 154,  30, 154,  29, 154,  28, 154,  27, 154,  26, 154,  25, 154,  24, 154,  23, 154,  22, 154,  21, 154,  20, 154,  19, 154,  18, 154,  17, 154,  16, 154,  15, 154,  14, 154,  13, 154,  12, 154,  11, 154,  10, 154,   9, 154,   8, 154,   7, 154,   6, 154,   5, 154,   4, 154,   3, 154,   2, 154,   1, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 250,  31, 250,  30, 250,  29, 250,  28, 250,  27, 250,  26, 250,  25, 250,  24, 250,  23, 250,  22, 242,  31, 242,  30, 242,  29, 242,  28, 242,  27, 242,  26, 242,  25, 242,  24, 242,  23, 242,  22, 242,  21, 242,  20, 242,  19, 242,  18, 242,  17, 242,  16, 242,  15, 242,  14, 242,  13, 242,  12, 242,  11, 242,  10, 242,   9, 242,   8, 242,   7, 242,   6, 242,   5, 242,   4, 242,   3, 242,   2, 242,   1, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 243,  31, 243,  30, 243,  29, 243,  28, 243,  27, 243,  26, 243,  25, 243,  24, 243,  23, 243,  22, 243,  21, 243,  20, 243,  19, 243,  18, 243,  17, 243,  16, 243,  15, 243,  14, 243,  13, 243,  12, 243,  11, 243,  10, 243,   9, 243,   8, 243,   7, 243,   6, 243,   5, 243,   4, 243,   3, 243,   2, 243,   1, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 175,  31, 175,  30, 175,  29, 175,  28, 175,  27, 175,  26, 175,  25, 175,  24, 175,  23, 175,  22, 175,  21, 175,  20, 175,  19, 175,  18, 175,  17, 175,  16, 175,  15, 175,  14, 175,  13, 175,  12, 210,  31, 210,  30, 210,  29, 210,  28, 210,  27, 210,  26, 210,  25, 210,  24, 210,  23, 210,  22, 210,  21, 210,  20, 210,  19, 210,  18, 210,  17, 210,  16, 210,  15, 210,  14, 210,  13, 210,  12, 210,  11, 210,  10, 210,   9, 210,   8, 210,   7, 210,   6, 210,   5, 210,   4, 210,   3, 210,   2, 210,   1, 210,   0, 210,   0, 210,   0, 210,   0, 210,   0, 210,   0, 210,   0, 210,   0, 210,   0, 210,   0, 210,   0, 210,   0, 210,   0, 210,   0, 210,   0, 210,   0, 210,   0, 210,   0, 210,   0, 210,   0, 210,   0, 210,   0, 210,   0, 210,   0, 103,  31, 103,  30, 103,  29, 103,  28, 103,  27, 103,  26, 103,  25, 103,  24, 103,  23, 103,  22, 103,  21, 103,  20, 103,  19, 103,  18, 103,  17, 103,  16, 103,  15, 103,  14, 103,  13, 103,  12, 103,  11, 103,  10, 103,   9, 103,   8, 103,   7, 103,   6, 103,   5, 103,   4, 103,   3, 103,   2, 103,   1, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0, 103,   0,   5,  31,   5,  30,   5,  29,   5,  28,   5,  27,   5,  26,   5,  25,   5,  24,   5,  23,   5,  22,   5,  21,   5,  20,   5,  19,   5,  18,   5,  17,   5,  16,   5,  15,   5,  14,   5,  13,   5,  12,   5,  11,   5,  10,   5,   9,   5,   8,   5,   7,   5,   6,   5,   5,   5,   4,   5,   3,   5,   2,   5,   1,   5,   0,   5,   0,   5,   0,   5,   0,   5,   0);
	constant SCENARIO_ADDRESS_19 : integer := 38947;


	--Scenario 20
	constant SCENARIO_LENGTH_20 : integer := 1015;
	type scenario_type_20 is array (0 to SCENARIO_LENGTH_20*2-1) of integer;
	signal scenario_input_20 : scenario_type_20 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 125,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 173,   0,   0,   0,   0,   0,   0,   0,  51,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  22,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  31,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 241,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  51,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 154,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 253,   0,   0,   0,  87,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 155,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  36,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 240,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 158,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 195,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 133,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  65,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 198,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 148,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 150,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 179,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 147,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  85,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  91,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  99,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 213,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 232,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  73,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  65,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 108,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_20  : scenario_type_20 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 125,  31, 125,  30, 125,  29, 125,  28, 125,  27, 125,  26, 125,  25, 125,  24, 125,  23, 125,  22, 125,  21, 125,  20, 125,  19, 125,  18, 125,  17, 125,  16, 125,  15, 125,  14, 125,  13, 125,  12, 125,  11, 125,  10, 125,   9, 125,   8, 125,   7, 125,   6, 125,   5, 125,   4, 125,   3, 125,   2, 125,   1, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 173,  31, 173,  30, 173,  29, 173,  28,  51,  31,  51,  30,  51,  29,  51,  28,  51,  27,  51,  26,  51,  25,  51,  24,  51,  23,  51,  22,  51,  21,  51,  20,  51,  19,  51,  18,  51,  17,  51,  16,  51,  15,  51,  14,  51,  13,  51,  12,  51,  11,  51,  10,  51,   9,  51,   8,  51,   7,  51,   6,  51,   5,  51,   4,  51,   3,  51,   2,  51,   1,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  22,  31,  22,  30,  22,  29,  22,  28,  22,  27,  22,  26,  22,  25,  22,  24,  22,  23,  22,  22,  22,  21,  22,  20,  22,  19,  22,  18,  22,  17,  22,  16,  22,  15,  22,  14,  22,  13,  22,  12,  22,  11,  22,  10,  22,   9,  22,   8,  22,   7,  22,   6,  22,   5,  22,   4,  22,   3,  22,   2,  22,   1,  22,   0,  22,   0,  22,   0,  31,  31,  31,  30,  31,  29,  31,  28,  31,  27,  31,  26,  31,  25,  31,  24,  31,  23,  31,  22,  31,  21,  31,  20,  31,  19,  31,  18,  31,  17,  31,  16,  31,  15,  31,  14,  31,  13,  31,  12,  31,  11,  31,  10,  31,   9,  31,   8,  31,   7,  31,   6, 241,  31, 241,  30, 241,  29, 241,  28, 241,  27, 241,  26, 241,  25, 241,  24, 241,  23, 241,  22, 241,  21, 241,  20, 241,  19, 241,  18, 241,  17, 241,  16, 241,  15, 241,  14, 241,  13, 241,  12, 241,  11, 241,  10, 241,   9, 241,   8, 241,   7, 241,   6, 241,   5, 241,   4, 241,   3, 241,   2, 241,   1, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0, 241,   0,  51,  31,  51,  30,  51,  29,  51,  28,  51,  27,  51,  26,  51,  25,  51,  24,  51,  23,  51,  22,  51,  21,  51,  20,  51,  19,  51,  18,  51,  17,  51,  16,  51,  15,  51,  14,  51,  13,  51,  12,  51,  11,  51,  10,  51,   9,  51,   8,  51,   7,  51,   6,  51,   5,  51,   4,  51,   3,  51,   2,  51,   1,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0,  51,   0, 154,  31, 154,  30, 154,  29, 154,  28, 154,  27, 154,  26, 154,  25, 154,  24, 154,  23, 154,  22, 154,  21, 154,  20, 154,  19, 154,  18, 154,  17, 154,  16, 154,  15, 154,  14, 154,  13, 154,  12, 154,  11, 154,  10, 154,   9, 154,   8, 154,   7, 154,   6, 154,   5, 154,   4, 154,   3, 154,   2, 154,   1, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 154,   0, 253,  31, 253,  30,  87,  31,  87,  30,  87,  29,  87,  28,  87,  27,  87,  26,  87,  25,  87,  24,  87,  23,  87,  22,  87,  21,  87,  20,  87,  19,  87,  18,  87,  17,  87,  16,  87,  15,  87,  14,  87,  13,  87,  12,  87,  11,  87,  10,  87,   9,  87,   8,  87,   7,  87,   6,  87,   5,  87,   4,  87,   3,  87,   2,  87,   1,  87,   0,  87,   0,  87,   0, 155,  31, 155,  30, 155,  29, 155,  28, 155,  27, 155,  26, 155,  25, 155,  24, 155,  23, 155,  22, 155,  21, 155,  20, 155,  19, 155,  18, 155,  17, 155,  16, 155,  15, 155,  14, 155,  13, 155,  12, 155,  11, 155,  10, 155,   9, 155,   8, 155,   7, 155,   6, 155,   5, 155,   4, 155,   3, 155,   2, 155,   1, 155,   0, 155,   0, 155,   0, 155,   0, 155,   0, 155,   0, 155,   0, 155,   0, 155,   0, 155,   0, 155,   0, 155,   0, 155,   0, 155,   0, 155,   0, 155,   0, 155,   0, 155,   0,  36,  31,  36,  30,  36,  29,  36,  28,  36,  27,  36,  26,  36,  25,  36,  24,  36,  23,  36,  22,  36,  21,  36,  20,  36,  19,  36,  18,  36,  17,  36,  16,  36,  15,  36,  14,  36,  13,  36,  12,  36,  11,  36,  10,  36,   9,  36,   8,  36,   7,  36,   6,  36,   5,  36,   4,  36,   3,  36,   2,  36,   1,  36,   0,  36,   0,  36,   0,  36,   0,  36,   0,  36,   0,  36,   0,  36,   0,  36,   0,  36,   0,  36,   0,  36,   0,  36,   0,  36,   0,  36,   0, 240,  31, 240,  30, 240,  29, 240,  28, 240,  27, 240,  26, 240,  25, 240,  24, 240,  23, 240,  22, 240,  21, 240,  20, 240,  19, 240,  18, 240,  17, 240,  16, 240,  15, 240,  14, 240,  13, 240,  12, 240,  11, 240,  10, 240,   9, 240,   8, 240,   7, 240,   6, 240,   5, 240,   4, 240,   3, 240,   2, 240,   1, 240,   0, 240,   0, 240,   0, 240,   0, 240,   0, 240,   0, 240,   0, 240,   0, 240,   0, 240,   0, 240,   0, 158,  31, 158,  30, 158,  29, 158,  28, 158,  27, 158,  26, 158,  25, 158,  24, 158,  23, 158,  22, 158,  21, 158,  20, 158,  19, 158,  18, 158,  17, 158,  16, 158,  15, 158,  14, 158,  13, 158,  12, 158,  11, 158,  10, 158,   9, 158,   8, 158,   7, 158,   6, 158,   5, 158,   4, 158,   3, 158,   2, 158,   1, 158,   0, 195,  31, 195,  30, 195,  29, 195,  28, 195,  27, 195,  26, 195,  25, 195,  24, 195,  23, 195,  22, 195,  21, 195,  20, 195,  19, 195,  18, 195,  17, 195,  16, 195,  15, 195,  14, 195,  13, 195,  12, 195,  11, 195,  10, 195,   9, 195,   8, 195,   7, 195,   6, 195,   5, 195,   4, 133,  31, 133,  30, 133,  29, 133,  28, 133,  27, 133,  26, 133,  25, 133,  24, 133,  23, 133,  22, 133,  21, 133,  20, 133,  19, 133,  18, 133,  17, 133,  16, 133,  15, 133,  14, 133,  13, 133,  12, 133,  11, 133,  10, 133,   9, 133,   8, 133,   7, 133,   6, 133,   5, 133,   4,  65,  31,  65,  30,  65,  29,  65,  28,  65,  27,  65,  26,  65,  25,  65,  24,  65,  23,  65,  22,  65,  21,  65,  20,  65,  19,  65,  18,  65,  17,  65,  16,  65,  15,  65,  14,  65,  13,  65,  12,  65,  11,  65,  10,  65,   9,  65,   8,  65,   7,  65,   6,  65,   5,  65,   4,  65,   3,  65,   2,  65,   1,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0,  65,   0, 198,  31, 198,  30, 198,  29, 198,  28, 198,  27, 198,  26, 198,  25, 198,  24, 198,  23, 198,  22, 198,  21, 198,  20, 198,  19, 198,  18, 198,  17, 198,  16, 198,  15, 198,  14, 198,  13, 198,  12, 198,  11, 198,  10, 198,   9, 198,   8, 148,  31, 148,  30, 148,  29, 148,  28, 148,  27, 148,  26, 148,  25, 148,  24, 148,  23, 148,  22, 148,  21, 148,  20, 148,  19, 148,  18, 150,  31, 150,  30, 150,  29, 150,  28, 150,  27, 150,  26, 150,  25, 150,  24, 150,  23, 150,  22, 150,  21, 150,  20, 150,  19, 150,  18, 150,  17, 150,  16, 150,  15, 150,  14, 150,  13, 150,  12, 150,  11, 150,  10, 150,   9, 150,   8, 150,   7, 150,   6, 150,   5, 150,   4, 150,   3, 150,   2, 150,   1, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 179,  31, 179,  30, 179,  29, 179,  28, 179,  27, 179,  26, 179,  25, 179,  24, 179,  23, 179,  22, 179,  21, 179,  20, 179,  19, 179,  18, 179,  17, 179,  16, 179,  15, 179,  14, 179,  13, 179,  12, 179,  11, 179,  10, 179,   9, 179,   8, 179,   7, 179,   6, 179,   5, 179,   4, 179,   3, 179,   2, 179,   1, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 147,  31, 147,  30, 147,  29, 147,  28, 147,  27, 147,  26, 147,  25, 147,  24, 147,  23, 147,  22, 147,  21, 147,  20, 147,  19, 147,  18, 147,  17, 147,  16, 147,  15, 147,  14, 147,  13, 147,  12, 147,  11, 147,  10, 147,   9, 147,   8, 147,   7, 147,   6, 147,   5, 147,   4, 147,   3, 147,   2, 147,   1, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0, 147,   0,  85,  31,  85,  30,  85,  29,  85,  28,  85,  27,  85,  26,  85,  25,  85,  24,  85,  23,  85,  22,  85,  21,  85,  20,  85,  19,  85,  18,  91,  31,  91,  30,  91,  29,  91,  28,  91,  27,  91,  26,  91,  25,  91,  24,  91,  23,  91,  22,  91,  21,  91,  20,  91,  19,  91,  18,  91,  17,  91,  16,  91,  15,  91,  14,  91,  13,  91,  12,  91,  11,  91,  10,  91,   9,  91,   8,  91,   7,  91,   6,  91,   5,  91,   4,  91,   3,  91,   2,  91,   1,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  99,  31,  99,  30,  99,  29,  99,  28,  99,  27,  99,  26,  99,  25,  99,  24,  99,  23,  99,  22,  99,  21,  99,  20,  99,  19,  99,  18,  99,  17,  99,  16,  99,  15,  99,  14,  99,  13,  99,  12,  99,  11,  99,  10,  99,   9, 213,  31, 213,  30, 213,  29, 213,  28, 213,  27, 213,  26, 213,  25, 213,  24, 213,  23, 213,  22, 213,  21, 213,  20, 213,  19, 213,  18, 213,  17, 213,  16, 213,  15, 213,  14, 213,  13, 213,  12, 213,  11, 213,  10, 213,   9, 213,   8, 213,   7, 213,   6, 213,   5, 213,   4, 213,   3, 213,   2, 213,   1, 213,   0, 213,   0, 213,   0, 213,   0, 213,   0, 213,   0, 213,   0, 213,   0, 213,   0, 213,   0, 213,   0, 213,   0, 213,   0, 232,  31, 232,  30, 232,  29, 232,  28, 232,  27, 232,  26, 232,  25, 232,  24, 232,  23, 232,  22, 232,  21,  73,  31,  73,  30,  73,  29,  73,  28,  73,  27,  73,  26,  73,  25,  73,  24,  73,  23,  73,  22,  73,  21,  73,  20,  65,  31,  65,  30,  65,  29,  65,  28,  65,  27,  65,  26,  65,  25,  65,  24,  65,  23,  65,  22,  65,  21,  65,  20,  65,  19,  65,  18,  65,  17,  65,  16,  65,  15,  65,  14,  65,  13,  65,  12,  65,  11,  65,  10,  65,   9,  65,   8,  65,   7,  65,   6,  65,   5, 108,  31, 108,  30, 108,  29, 108,  28, 108,  27, 108,  26, 108,  25, 108,  24, 108,  23, 108,  22, 108,  21);
	constant SCENARIO_ADDRESS_20 : integer := 40962;


	--Scenario 21
	constant SCENARIO_LENGTH_21 : integer := 1022;
	type scenario_type_21 is array (0 to SCENARIO_LENGTH_21*2-1) of integer;
	signal scenario_input_21 : scenario_type_21 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 200,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  78,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 196,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  99,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 108,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  33,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  79,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  21,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  43,   0,   0,   0, 149,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 248,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 126,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 158,   0,   0,   0,   0,   0,   0,   0, 157,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 219,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 251,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  16,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  19,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 194,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 167,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  50,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 129,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 118,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 117,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   7,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 160,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 175,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 135,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 130,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_21  : scenario_type_21 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 200,  31, 200,  30, 200,  29, 200,  28, 200,  27, 200,  26,  78,  31,  78,  30,  78,  29,  78,  28,  78,  27,  78,  26,  78,  25,  78,  24,  78,  23,  78,  22,  78,  21,  78,  20,  78,  19,  78,  18,  78,  17,  78,  16,  78,  15,  78,  14,  78,  13,  78,  12,  78,  11,  78,  10,  78,   9,  78,   8,  78,   7,  78,   6,  78,   5,  78,   4,  78,   3,  78,   2,  78,   1,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0,  78,   0, 196,  31, 196,  30, 196,  29, 196,  28, 196,  27, 196,  26, 196,  25, 196,  24, 196,  23, 196,  22, 196,  21, 196,  20, 196,  19,  99,  31,  99,  30,  99,  29,  99,  28,  99,  27,  99,  26,  99,  25,  99,  24,  99,  23,  99,  22,  99,  21,  99,  20,  99,  19,  99,  18,  99,  17,  99,  16,  99,  15,  99,  14,  99,  13,  99,  12,  99,  11,  99,  10,  99,   9,  99,   8,  99,   7,  99,   6,  99,   5,  99,   4,  99,   3,  99,   2,  99,   1,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0, 108,  31, 108,  30, 108,  29, 108,  28, 108,  27, 108,  26, 108,  25, 108,  24, 108,  23, 108,  22, 108,  21, 108,  20, 108,  19, 108,  18, 108,  17, 108,  16, 108,  15, 108,  14, 108,  13, 108,  12, 108,  11, 108,  10, 108,   9, 108,   8, 108,   7, 108,   6, 108,   5, 108,   4,  33,  31,  33,  30,  33,  29,  33,  28,  33,  27,  33,  26,  33,  25,  33,  24,  33,  23,  33,  22,  33,  21,  33,  20,  33,  19,  33,  18,  33,  17,  33,  16,  33,  15,  33,  14,  33,  13,  33,  12,  33,  11,  33,  10,  33,   9,  33,   8,  33,   7,  33,   6,  33,   5,  33,   4,  33,   3,  33,   2,  33,   1,  33,   0,  33,   0,  33,   0,  33,   0,  33,   0,  33,   0,  79,  31,  79,  30,  79,  29,  79,  28,  79,  27,  79,  26,  79,  25,  79,  24,  79,  23,  79,  22,  79,  21,  79,  20,  79,  19,  79,  18,  79,  17,  79,  16,  79,  15,  79,  14,  79,  13,  79,  12,  79,  11,  21,  31,  21,  30,  21,  29,  21,  28,  21,  27,  21,  26,  21,  25,  21,  24,  21,  23,  21,  22,  21,  21,  21,  20,  21,  19,  21,  18,  21,  17,  21,  16,  21,  15,  21,  14,  21,  13,  21,  12,  21,  11,  21,  10,  21,   9,  21,   8,  21,   7,  43,  31,  43,  30, 149,  31, 149,  30, 149,  29, 149,  28, 149,  27, 149,  26, 149,  25, 149,  24, 149,  23, 149,  22, 149,  21, 149,  20, 149,  19, 149,  18, 149,  17, 149,  16, 149,  15, 149,  14, 149,  13, 149,  12, 149,  11, 149,  10, 149,   9, 149,   8, 149,   7, 149,   6, 149,   5, 149,   4, 149,   3, 149,   2, 149,   1, 149,   0, 149,   0, 149,   0, 149,   0, 149,   0, 248,  31, 248,  30, 248,  29, 248,  28, 248,  27, 248,  26, 248,  25, 248,  24, 248,  23, 248,  22, 248,  21, 126,  31, 126,  30, 126,  29, 126,  28, 126,  27, 126,  26, 126,  25, 126,  24, 126,  23, 126,  22, 126,  21, 126,  20, 126,  19, 126,  18, 126,  17, 126,  16, 126,  15, 126,  14, 126,  13, 126,  12, 126,  11, 126,  10, 126,   9, 126,   8, 126,   7, 126,   6, 126,   5, 126,   4, 126,   3, 126,   2, 126,   1, 126,   0, 126,   0, 126,   0, 158,  31, 158,  30, 158,  29, 158,  28, 157,  31, 157,  30, 157,  29, 157,  28, 157,  27, 157,  26, 157,  25, 157,  24, 157,  23, 157,  22, 157,  21, 157,  20, 157,  19, 157,  18, 157,  17, 157,  16, 157,  15, 157,  14, 157,  13, 157,  12, 157,  11, 157,  10, 157,   9, 157,   8, 157,   7, 157,   6, 157,   5, 157,   4, 157,   3, 157,   2, 157,   1, 157,   0, 157,   0, 157,   0, 157,   0, 157,   0, 157,   0, 157,   0, 157,   0, 157,   0, 157,   0, 157,   0, 157,   0, 157,   0, 157,   0, 157,   0, 157,   0, 157,   0, 157,   0, 157,   0, 157,   0, 157,   0, 219,  31, 219,  30, 219,  29, 219,  28, 219,  27, 219,  26, 219,  25, 219,  24, 219,  23, 219,  22, 219,  21, 219,  20, 219,  19, 219,  18, 219,  17, 219,  16, 219,  15, 219,  14, 219,  13, 219,  12, 219,  11, 219,  10, 219,   9, 219,   8, 219,   7, 219,   6, 219,   5, 219,   4, 219,   3, 219,   2, 219,   1, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 251,  31, 251,  30, 251,  29, 251,  28, 251,  27, 251,  26, 251,  25, 251,  24, 251,  23, 251,  22, 251,  21, 251,  20, 251,  19, 251,  18, 251,  17, 251,  16, 251,  15, 251,  14, 251,  13, 251,  12, 251,  11, 251,  10, 251,   9, 251,   8, 251,   7, 251,   6, 251,   5, 251,   4, 251,   3, 251,   2,  16,  31,  16,  30,  16,  29,  16,  28,  16,  27,  16,  26,  16,  25,  16,  24,  16,  23,  16,  22,  16,  21,  19,  31,  19,  30,  19,  29,  19,  28,  19,  27,  19,  26,  19,  25,  19,  24,  19,  23,  19,  22,  19,  21,  19,  20,  19,  19,  19,  18,  19,  17,  19,  16,  19,  15,  19,  14,  19,  13,  19,  12,  19,  11,  19,  10,  19,   9,  19,   8,  19,   7, 194,  31, 194,  30, 194,  29, 194,  28, 194,  27, 194,  26, 194,  25, 194,  24, 167,  31, 167,  30, 167,  29, 167,  28, 167,  27, 167,  26, 167,  25, 167,  24, 167,  23, 167,  22, 167,  21, 167,  20, 167,  19, 167,  18, 167,  17, 167,  16, 167,  15, 167,  14, 167,  13, 167,  12, 167,  11, 167,  10, 167,   9, 167,   8, 167,   7,  50,  31,  50,  30,  50,  29,  50,  28,  50,  27,  50,  26,  50,  25,  50,  24,  50,  23,  50,  22,  50,  21,  50,  20,  50,  19,  50,  18,  50,  17,  50,  16,  50,  15,  50,  14,  50,  13,  50,  12,  50,  11,  50,  10,  50,   9,  50,   8, 129,  31, 129,  30, 129,  29, 129,  28, 129,  27, 129,  26, 129,  25, 129,  24, 129,  23, 129,  22, 129,  21, 129,  20, 129,  19, 129,  18, 129,  17, 129,  16, 129,  15, 129,  14, 129,  13, 129,  12, 129,  11, 129,  10, 129,   9, 129,   8, 129,   7, 129,   6, 129,   5, 129,   4, 129,   3, 129,   2, 129,   1, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 118,  31, 118,  30, 118,  29, 118,  28, 118,  27, 118,  26, 118,  25, 118,  24, 118,  23, 118,  22, 118,  21, 118,  20, 118,  19, 118,  18, 118,  17, 118,  16, 117,  31, 117,  30, 117,  29, 117,  28, 117,  27, 117,  26, 117,  25, 117,  24, 117,  23, 117,  22, 117,  21, 117,  20,   7,  31,   7,  30,   7,  29,   7,  28,   7,  27,   7,  26,   7,  25,   7,  24,   7,  23,   7,  22,   7,  21,   7,  20,   7,  19,   7,  18,   7,  17,   7,  16,   7,  15,   7,  14,   7,  13,   7,  12,   7,  11,   7,  10,   7,   9,   7,   8,   7,   7,   7,   6,   7,   5,   7,   4,   7,   3,   7,   2,   7,   1,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0,   7,   0, 160,  31, 160,  30, 160,  29, 160,  28, 160,  27, 160,  26, 160,  25, 160,  24, 160,  23, 160,  22, 160,  21, 160,  20, 160,  19, 160,  18, 160,  17, 160,  16, 160,  15, 160,  14, 160,  13, 160,  12, 160,  11, 160,  10, 160,   9, 160,   8, 160,   7, 160,   6, 160,   5, 160,   4, 160,   3, 160,   2, 160,   1, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 160,   0, 175,  31, 175,  30, 175,  29, 175,  28, 175,  27, 175,  26, 175,  25, 175,  24, 175,  23, 175,  22, 175,  21, 175,  20, 175,  19, 175,  18, 175,  17, 175,  16, 175,  15, 175,  14, 175,  13, 175,  12, 175,  11, 175,  10, 175,   9, 175,   8, 175,   7, 175,   6, 175,   5, 175,   4, 175,   3, 175,   2, 175,   1, 175,   0, 175,   0, 175,   0, 135,  31, 135,  30, 135,  29, 135,  28, 135,  27, 135,  26, 135,  25, 135,  24, 135,  23, 135,  22, 135,  21, 135,  20, 135,  19, 135,  18, 135,  17, 135,  16, 135,  15, 135,  14, 135,  13, 135,  12, 135,  11, 135,  10, 135,   9, 135,   8, 135,   7, 135,   6, 135,   5, 135,   4, 135,   3, 135,   2, 135,   1, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 135,   0, 130,  31, 130,  30, 130,  29, 130,  28, 130,  27, 130,  26, 130,  25, 130,  24, 130,  23, 130,  22, 130,  21, 130,  20, 130,  19, 130,  18, 130,  17, 130,  16, 130,  15, 130,  14, 130,  13, 130,  12, 130,  11, 130,  10, 130,   9, 130,   8, 130,   7, 130,   6, 130,   5, 130,   4, 130,   3, 130,   2, 130,   1, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0, 130,   0);
	constant SCENARIO_ADDRESS_21 : integer := 43012;


	--Scenario 22
	constant SCENARIO_LENGTH_22 : integer := 1009;
	type scenario_type_22 is array (0 to SCENARIO_LENGTH_22*2-1) of integer;
	signal scenario_input_22 : scenario_type_22 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  11,   0, 200,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   9,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  64,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 251,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 227,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 179,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 124,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  13,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 244,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 152,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  32,   0, 159,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  68,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 201,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 137,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 220,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   3,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 214,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  20,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 146,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  87,   0,   0,   0,   0,   0,  14,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 167,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 138,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  27,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_22  : scenario_type_22 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  11,  31, 200,  31, 200,  30, 200,  29, 200,  28, 200,  27, 200,  26, 200,  25, 200,  24, 200,  23, 200,  22, 200,  21, 200,  20, 200,  19, 200,  18, 200,  17, 200,  16, 200,  15, 200,  14, 200,  13, 200,  12, 200,  11, 200,  10, 200,   9, 200,   8, 200,   7, 200,   6, 200,   5, 200,   4, 200,   3, 200,   2, 200,   1, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0,   9,  31,   9,  30,   9,  29,   9,  28,   9,  27,   9,  26,   9,  25,   9,  24,   9,  23,   9,  22,   9,  21,   9,  20,   9,  19,   9,  18,   9,  17,   9,  16,   9,  15,   9,  14,   9,  13,   9,  12,   9,  11,   9,  10,   9,   9,   9,   8,   9,   7,   9,   6,   9,   5,   9,   4,   9,   3,   9,   2,   9,   1,   9,   0,   9,   0,   9,   0,   9,   0,   9,   0,   9,   0,   9,   0,   9,   0,   9,   0,   9,   0,  64,  31,  64,  30,  64,  29,  64,  28,  64,  27,  64,  26,  64,  25,  64,  24,  64,  23,  64,  22,  64,  21,  64,  20,  64,  19,  64,  18,  64,  17, 251,  31, 251,  30, 251,  29, 251,  28, 251,  27, 251,  26, 251,  25, 251,  24, 251,  23, 251,  22, 251,  21, 251,  20, 251,  19, 251,  18, 251,  17, 251,  16, 251,  15, 251,  14, 251,  13, 251,  12, 251,  11, 251,  10, 251,   9, 251,   8, 251,   7, 251,   6, 251,   5, 251,   4, 251,   3, 251,   2, 251,   1, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 251,   0, 227,  31, 227,  30, 227,  29, 227,  28, 227,  27, 227,  26, 227,  25, 227,  24, 227,  23, 227,  22, 227,  21, 227,  20, 227,  19, 227,  18, 227,  17, 227,  16, 227,  15, 227,  14, 227,  13, 227,  12, 227,  11, 227,  10, 227,   9, 227,   8, 227,   7, 227,   6, 227,   5, 227,   4, 227,   3, 227,   2, 227,   1, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 227,   0, 179,  31, 179,  30, 179,  29, 179,  28, 179,  27, 179,  26, 179,  25, 179,  24, 179,  23, 179,  22, 179,  21, 179,  20, 179,  19, 179,  18, 179,  17, 179,  16, 179,  15, 179,  14, 179,  13, 179,  12, 179,  11, 179,  10, 179,   9, 179,   8, 179,   7, 179,   6, 179,   5, 179,   4, 179,   3, 179,   2, 179,   1, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 179,   0, 124,  31, 124,  30, 124,  29, 124,  28, 124,  27, 124,  26, 124,  25, 124,  24, 124,  23, 124,  22, 124,  21, 124,  20, 124,  19, 124,  18, 124,  17, 124,  16, 124,  15, 124,  14, 124,  13, 124,  12, 124,  11, 124,  10, 124,   9, 124,   8, 124,   7, 124,   6, 124,   5, 124,   4, 124,   3, 124,   2, 124,   1, 124,   0, 124,   0, 124,   0, 124,   0, 124,   0, 124,   0, 124,   0, 124,   0,  13,  31,  13,  30,  13,  29,  13,  28,  13,  27,  13,  26,  13,  25,  13,  24,  13,  23,  13,  22,  13,  21,  13,  20,  13,  19,  13,  18,  13,  17,  13,  16,  13,  15,  13,  14, 244,  31, 244,  30, 244,  29, 244,  28, 244,  27, 244,  26, 244,  25, 244,  24, 244,  23, 244,  22, 244,  21, 244,  20, 244,  19, 244,  18, 244,  17, 244,  16, 244,  15, 244,  14, 244,  13, 244,  12, 244,  11, 244,  10, 244,   9, 244,   8, 244,   7, 244,   6, 244,   5, 244,   4, 244,   3, 244,   2, 244,   1, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 244,   0, 152,  31, 152,  30, 152,  29, 152,  28, 152,  27, 152,  26, 152,  25, 152,  24, 152,  23, 152,  22, 152,  21, 152,  20, 152,  19, 152,  18, 152,  17, 152,  16, 152,  15, 152,  14, 152,  13, 152,  12, 152,  11, 152,  10, 152,   9, 152,   8, 152,   7,  32,  31, 159,  31, 159,  30, 159,  29, 159,  28, 159,  27, 159,  26, 159,  25, 159,  24, 159,  23, 159,  22, 159,  21, 159,  20, 159,  19,  68,  31,  68,  30,  68,  29,  68,  28,  68,  27,  68,  26,  68,  25,  68,  24,  68,  23,  68,  22,  68,  21,  68,  20,  68,  19,  68,  18,  68,  17,  68,  16,  68,  15,  68,  14,  68,  13,  68,  12,  68,  11,  68,  10,  68,   9,  68,   8,  68,   7,  68,   6,  68,   5,  68,   4,  68,   3,  68,   2,  68,   1,  68,   0, 201,  31, 201,  30, 201,  29, 201,  28, 201,  27, 201,  26, 201,  25, 201,  24, 201,  23, 201,  22, 201,  21, 201,  20, 201,  19, 201,  18, 201,  17, 201,  16, 201,  15, 201,  14, 201,  13, 201,  12, 201,  11, 201,  10, 201,   9, 201,   8, 201,   7, 201,   6, 201,   5, 201,   4, 201,   3, 201,   2, 201,   1, 201,   0, 201,   0, 201,   0, 201,   0, 201,   0, 201,   0, 201,   0, 201,   0, 201,   0, 201,   0, 201,   0, 201,   0, 201,   0, 201,   0, 137,  31, 137,  30, 137,  29, 137,  28, 137,  27, 137,  26, 137,  25, 137,  24, 137,  23, 137,  22, 137,  21, 137,  20, 137,  19, 137,  18, 137,  17, 137,  16, 137,  15, 137,  14, 137,  13, 137,  12, 137,  11, 137,  10, 137,   9, 137,   8, 137,   7, 137,   6, 137,   5, 137,   4, 137,   3, 137,   2, 137,   1, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 137,   0, 220,  31, 220,  30, 220,  29, 220,  28, 220,  27, 220,  26, 220,  25, 220,  24, 220,  23, 220,  22, 220,  21, 220,  20, 220,  19, 220,  18, 220,  17, 220,  16, 220,  15, 220,  14, 220,  13, 220,  12, 220,  11, 220,  10, 220,   9, 220,   8, 220,   7, 220,   6, 220,   5, 220,   4, 220,   3, 220,   2, 220,   1, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0,   3,  31,   3,  30,   3,  29,   3,  28,   3,  27,   3,  26,   3,  25,   3,  24,   3,  23,   3,  22,   3,  21,   3,  20,   3,  19,   3,  18,   3,  17,   3,  16,   3,  15,   3,  14,   3,  13,   3,  12,   3,  11,   3,  10,   3,   9,   3,   8,   3,   7,   3,   6,   3,   5,   3,   4,   3,   3,   3,   2,   3,   1,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0,   3,   0, 214,  31, 214,  30, 214,  29, 214,  28, 214,  27, 214,  26, 214,  25, 214,  24, 214,  23, 214,  22, 214,  21, 214,  20, 214,  19, 214,  18, 214,  17, 214,  16, 214,  15, 214,  14, 214,  13, 214,  12, 214,  11, 214,  10, 214,   9, 214,   8, 214,   7, 214,   6, 214,   5, 214,   4, 214,   3, 214,   2, 214,   1, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0, 214,   0,  20,  31,  20,  30,  20,  29,  20,  28,  20,  27,  20,  26,  20,  25,  20,  24,  20,  23,  20,  22,  20,  21,  20,  20,  20,  19,  20,  18,  20,  17,  20,  16,  20,  15,  20,  14,  20,  13,  20,  12,  20,  11,  20,  10,  20,   9,  20,   8,  20,   7,  20,   6,  20,   5,  20,   4,  20,   3,  20,   2,  20,   1,  20,   0,  20,   0,  20,   0,  20,   0,  20,   0, 146,  31, 146,  30, 146,  29, 146,  28, 146,  27, 146,  26, 146,  25, 146,  24, 146,  23, 146,  22, 146,  21, 146,  20, 146,  19, 146,  18, 146,  17, 146,  16, 146,  15, 146,  14, 146,  13, 146,  12, 146,  11, 146,  10, 146,   9, 146,   8, 146,   7, 146,   6, 146,   5, 146,   4, 146,   3, 146,   2, 146,   1, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0,  87,  31,  87,  30,  87,  29,  14,  31,  14,  30,  14,  29,  14,  28,  14,  27,  14,  26,  14,  25,  14,  24,  14,  23,  14,  22,  14,  21,  14,  20,  14,  19,  14,  18,  14,  17,  14,  16,  14,  15,  14,  14,  14,  13,  14,  12,  14,  11,  14,  10,  14,   9,  14,   8,  14,   7,  14,   6,  14,   5,  14,   4,  14,   3,  14,   2,  14,   1,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0, 167,  31, 167,  30, 167,  29, 167,  28, 167,  27, 167,  26, 167,  25, 167,  24, 167,  23, 167,  22, 167,  21, 167,  20, 167,  19, 167,  18, 167,  17, 167,  16, 167,  15, 167,  14, 167,  13, 167,  12, 167,  11, 167,  10, 167,   9, 167,   8, 167,   7, 167,   6, 167,   5, 167,   4, 167,   3, 167,   2, 167,   1, 167,   0, 167,   0, 167,   0, 167,   0, 167,   0, 167,   0, 167,   0, 167,   0, 167,   0, 167,   0, 167,   0, 167,   0, 138,  31, 138,  30, 138,  29, 138,  28, 138,  27, 138,  26, 138,  25, 138,  24, 138,  23, 138,  22, 138,  21, 138,  20, 138,  19, 138,  18, 138,  17, 138,  16, 138,  15, 138,  14, 138,  13, 138,  12, 138,  11, 138,  10, 138,   9, 138,   8, 138,   7, 138,   6, 138,   5, 138,   4,  27,  31,  27,  30,  27,  29,  27,  28,  27,  27,  27,  26,  27,  25,  27,  24,  27,  23,  27,  22,  27,  21,  27,  20,  27,  19,  27,  18,  27,  17,  27,  16,  27,  15,  27,  14,  27,  13,  27,  12,  27,  11,  27,  10,  27,   9,  27,   8,  27,   7,  27,   6,  27,   5,  27,   4,  27,   3,  27,   2,  27,   1,  27,   0,  27,   0,  27,   0,  27,   0,  27,   0,  27,   0,  27,   0,  27,   0);
	constant SCENARIO_ADDRESS_22 : integer := 45065;


	--Scenario 23
	constant SCENARIO_LENGTH_23 : integer := 1;
	type scenario_type_23 is array (0 to SCENARIO_LENGTH_23*2-1) of integer;
	signal scenario_input_23 : scenario_type_23 := (7,   7);
	signal scenario_full_23  : scenario_type_23 := (7,   7);
	constant SCENARIO_ADDRESS_23 : integer := 48928;
	--This sequence is going to be ignored by the component
	--as the i_k parameter is will be set to zero


	--Scenario 24
	constant SCENARIO_LENGTH_24 : integer := 974;
	type scenario_type_24 is array (0 to SCENARIO_LENGTH_24*2-1) of integer;
	signal scenario_input_24 : scenario_type_24 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  67,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 154,   0,   0,   0,  98,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 104,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  67,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 246,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 207,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  77,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  73,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 142,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 122,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  32,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 144,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  10,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  23,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  40,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 212,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  69,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 150,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  88,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 203,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 237,   0,   0,   0,  80,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  81,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_24  : scenario_type_24 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  67,  31,  67,  30,  67,  29,  67,  28,  67,  27,  67,  26,  67,  25,  67,  24,  67,  23,  67,  22,  67,  21,  67,  20,  67,  19,  67,  18,  67,  17,  67,  16,  67,  15,  67,  14,  67,  13,  67,  12,  67,  11,  67,  10,  67,   9,  67,   8,  67,   7,  67,   6,  67,   5,  67,   4,  67,   3,  67,   2,  67,   1,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0, 154,  31, 154,  30,  98,  31,  98,  30,  98,  29,  98,  28,  98,  27,  98,  26,  98,  25,  98,  24,  98,  23, 104,  31, 104,  30, 104,  29, 104,  28, 104,  27, 104,  26, 104,  25, 104,  24, 104,  23, 104,  22, 104,  21, 104,  20, 104,  19, 104,  18, 104,  17, 104,  16, 104,  15, 104,  14, 104,  13, 104,  12, 104,  11, 104,  10, 104,   9, 104,   8, 104,   7, 104,   6, 104,   5, 104,   4, 104,   3,  67,  31,  67,  30,  67,  29,  67,  28,  67,  27,  67,  26,  67,  25,  67,  24,  67,  23,  67,  22,  67,  21,  67,  20,  67,  19,  67,  18,  67,  17,  67,  16,  67,  15,  67,  14,  67,  13,  67,  12,  67,  11,  67,  10,  67,   9,  67,   8,  67,   7,  67,   6,  67,   5,  67,   4,  67,   3,  67,   2,  67,   1,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0, 246,  31, 246,  30, 246,  29, 246,  28, 246,  27, 246,  26, 246,  25, 246,  24, 246,  23, 246,  22, 246,  21, 246,  20, 246,  19, 246,  18, 246,  17, 246,  16, 246,  15, 246,  14, 246,  13, 246,  12, 246,  11, 246,  10, 246,   9, 246,   8, 246,   7, 246,   6, 246,   5, 246,   4, 246,   3, 246,   2, 207,  31, 207,  30, 207,  29, 207,  28, 207,  27, 207,  26, 207,  25, 207,  24, 207,  23, 207,  22, 207,  21, 207,  20, 207,  19, 207,  18, 207,  17, 207,  16, 207,  15, 207,  14, 207,  13, 207,  12, 207,  11, 207,  10, 207,   9, 207,   8,  77,  31,  77,  30,  77,  29,  77,  28,  77,  27,  77,  26,  77,  25,  77,  24,  77,  23,  77,  22,  77,  21,  77,  20,  77,  19,  77,  18,  77,  17,  77,  16,  77,  15,  77,  14,  77,  13,  77,  12,  77,  11,  77,  10,  77,   9,  77,   8,  77,   7,  77,   6,  77,   5,  77,   4,  77,   3,  73,  31,  73,  30,  73,  29,  73,  28,  73,  27,  73,  26,  73,  25,  73,  24,  73,  23,  73,  22,  73,  21,  73,  20,  73,  19,  73,  18,  73,  17,  73,  16,  73,  15,  73,  14,  73,  13,  73,  12,  73,  11,  73,  10,  73,   9,  73,   8,  73,   7,  73,   6,  73,   5,  73,   4,  73,   3,  73,   2,  73,   1,  73,   0,  73,   0,  73,   0,  73,   0,  73,   0,  73,   0,  73,   0, 142,  31, 142,  30, 142,  29, 142,  28, 142,  27, 142,  26, 142,  25, 142,  24, 142,  23, 142,  22, 142,  21, 142,  20, 142,  19, 142,  18, 122,  31, 122,  30, 122,  29, 122,  28, 122,  27, 122,  26, 122,  25, 122,  24, 122,  23,  32,  31,  32,  30,  32,  29,  32,  28,  32,  27,  32,  26,  32,  25,  32,  24,  32,  23,  32,  22,  32,  21,  32,  20,  32,  19,  32,  18,  32,  17,  32,  16,  32,  15,  32,  14,  32,  13,  32,  12,  32,  11,  32,  10,  32,   9,  32,   8,  32,   7,  32,   6,  32,   5,  32,   4,  32,   3,  32,   2,  32,   1,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0, 144,  31, 144,  30, 144,  29, 144,  28, 144,  27, 144,  26, 144,  25, 144,  24, 144,  23, 144,  22, 144,  21, 144,  20, 144,  19, 144,  18, 144,  17, 144,  16, 144,  15, 144,  14, 144,  13, 144,  12, 144,  11, 144,  10, 144,   9, 144,   8, 144,   7,  10,  31,  10,  30,  10,  29,  10,  28,  10,  27,  10,  26,  10,  25,  10,  24,  10,  23,  10,  22,  10,  21,  10,  20,  10,  19,  10,  18,  10,  17,  10,  16,  10,  15,  10,  14,  10,  13,  10,  12,  10,  11,  10,  10,  10,   9,  10,   8,  10,   7,  10,   6,  10,   5,  10,   4,  10,   3,  10,   2,  10,   1,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  10,   0,  23,  31,  23,  30,  23,  29,  23,  28,  23,  27,  23,  26,  23,  25,  23,  24,  23,  23,  23,  22,  23,  21,  23,  20,  23,  19,  23,  18,  23,  17,  23,  16,  23,  15,  23,  14,  23,  13,  23,  12,  23,  11,  23,  10,  23,   9,  23,   8,  23,   7,  40,  31,  40,  30,  40,  29,  40,  28,  40,  27,  40,  26,  40,  25,  40,  24,  40,  23,  40,  22,  40,  21,  40,  20,  40,  19,  40,  18,  40,  17,  40,  16,  40,  15,  40,  14,  40,  13,  40,  12,  40,  11,  40,  10,  40,   9,  40,   8, 212,  31, 212,  30, 212,  29, 212,  28, 212,  27, 212,  26, 212,  25, 212,  24, 212,  23, 212,  22, 212,  21, 212,  20, 212,  19, 212,  18, 212,  17, 212,  16, 212,  15, 212,  14, 212,  13, 212,  12, 212,  11, 212,  10, 212,   9, 212,   8, 212,   7, 212,   6, 212,   5, 212,   4, 212,   3, 212,   2, 212,   1, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0, 212,   0,  69,  31,  69,  30,  69,  29,  69,  28,  69,  27,  69,  26,  69,  25,  69,  24,  69,  23,  69,  22,  69,  21,  69,  20,  69,  19,  69,  18,  69,  17,  69,  16,  69,  15,  69,  14,  69,  13,  69,  12,  69,  11,  69,  10,  69,   9,  69,   8,  69,   7,  69,   6,  69,   5,  69,   4,  69,   3,  69,   2,  69,   1,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0,  69,   0, 150,  31, 150,  30, 150,  29, 150,  28, 150,  27, 150,  26, 150,  25, 150,  24, 150,  23, 150,  22, 150,  21, 150,  20, 150,  19, 150,  18, 150,  17, 150,  16, 150,  15, 150,  14, 150,  13, 150,  12, 150,  11, 150,  10, 150,   9, 150,   8, 150,   7, 150,   6, 150,   5, 150,   4, 150,   3, 150,   2, 150,   1, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0, 150,   0,  88,  31,  88,  30,  88,  29,  88,  28,  88,  27,  88,  26,  88,  25,  88,  24,  88,  23,  88,  22,  88,  21,  88,  20,  88,  19,  88,  18,  88,  17,  88,  16,  88,  15, 203,  31, 203,  30, 203,  29, 203,  28, 203,  27, 203,  26, 203,  25, 203,  24, 203,  23, 203,  22, 203,  21, 203,  20, 203,  19, 203,  18, 203,  17, 203,  16, 203,  15, 237,  31, 237,  30,  80,  31,  80,  30,  80,  29,  80,  28,  80,  27,  80,  26,  80,  25,  80,  24,  80,  23,  80,  22,  80,  21,  80,  20,  80,  19,  80,  18,  80,  17,  80,  16,  80,  15,  80,  14,  80,  13,  80,  12,  80,  11,  80,  10,  80,   9,  80,   8,  80,   7,  80,   6,  80,   5,  80,   4,  80,   3,  80,   2,  80,   1,  80,   0,  80,   0,  80,   0,  80,   0,  80,   0,  80,   0,  80,   0,  80,   0,  80,   0,  80,   0,  80,   0,  80,   0,  80,   0,  80,   0,  80,   0,  80,   0,  80,   0,  80,   0,  80,   0,  81,  31,  81,  30,  81,  29,  81,  28,  81,  27,  81,  26,  81,  25,  81,  24,  81,  23,  81,  22,  81,  21,  81,  20,  81,  19,  81,  18,  81,  17,  81,  16,  81,  15,  81,  14,  81,  13,  81,  12,  81,  11,  81,  10,  81,   9,  81,   8,  81,   7,  81,   6,  81,   5,  81,   4,  81,   3,  81,   2,  81,   1,  81,   0);
	constant SCENARIO_ADDRESS_24 : integer := 49188;


	--Scenario 25
	constant SCENARIO_LENGTH_25 : integer := 989;
	type scenario_type_25 is array (0 to SCENARIO_LENGTH_25*2-1) of integer;
	signal scenario_input_25 : scenario_type_25 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 239,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 136,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   6,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 119,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 137,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 103,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  45,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 211,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 156,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 143,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 233,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 200,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  91,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  35,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  70,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 216,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 219,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 176,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 253,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 139,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 170,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 191,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 127,   0,   0,   0, 141,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  36,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  55,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 120,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 218,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  32,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_25  : scenario_type_25 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 239,  31, 239,  30, 239,  29, 239,  28, 239,  27, 239,  26, 239,  25, 239,  24, 239,  23, 239,  22, 239,  21, 239,  20, 239,  19, 239,  18, 239,  17, 239,  16, 136,  31, 136,  30, 136,  29, 136,  28, 136,  27, 136,  26, 136,  25, 136,  24, 136,  23, 136,  22, 136,  21, 136,  20, 136,  19, 136,  18, 136,  17, 136,  16, 136,  15, 136,  14, 136,  13, 136,  12, 136,  11,   6,  31,   6,  30,   6,  29,   6,  28,   6,  27,   6,  26,   6,  25,   6,  24,   6,  23,   6,  22,   6,  21,   6,  20,   6,  19,   6,  18,   6,  17,   6,  16,   6,  15,   6,  14,   6,  13,   6,  12,   6,  11,   6,  10,   6,   9,   6,   8,   6,   7,   6,   6,   6,   5,   6,   4,   6,   3,   6,   2,   6,   1,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0,   6,   0, 119,  31, 119,  30, 119,  29, 119,  28, 119,  27, 119,  26, 119,  25, 119,  24, 119,  23, 119,  22, 119,  21, 119,  20, 119,  19, 119,  18, 119,  17, 119,  16, 119,  15, 119,  14, 119,  13, 119,  12, 119,  11, 119,  10, 119,   9, 119,   8, 119,   7, 119,   6, 119,   5, 119,   4, 119,   3, 119,   2, 137,  31, 137,  30, 137,  29, 137,  28, 137,  27, 137,  26, 137,  25, 137,  24, 137,  23, 137,  22, 137,  21, 137,  20, 137,  19, 137,  18, 137,  17, 137,  16, 137,  15, 137,  14, 137,  13, 137,  12, 137,  11, 137,  10, 137,   9, 137,   8, 137,   7, 103,  31, 103,  30, 103,  29, 103,  28, 103,  27, 103,  26, 103,  25, 103,  24, 103,  23, 103,  22, 103,  21, 103,  20, 103,  19, 103,  18, 103,  17, 103,  16, 103,  15, 103,  14, 103,  13, 103,  12, 103,  11, 103,  10, 103,   9, 103,   8, 103,   7, 103,   6, 103,   5, 103,   4, 103,   3, 103,   2, 103,   1, 103,   0,  45,  31,  45,  30,  45,  29,  45,  28,  45,  27,  45,  26,  45,  25,  45,  24,  45,  23,  45,  22,  45,  21,  45,  20,  45,  19,  45,  18,  45,  17,  45,  16,  45,  15,  45,  14,  45,  13,  45,  12,  45,  11,  45,  10,  45,   9,  45,   8,  45,   7,  45,   6,  45,   5,  45,   4, 211,  31, 211,  30, 211,  29, 211,  28, 211,  27, 211,  26, 211,  25, 211,  24, 211,  23, 211,  22, 156,  31, 156,  30, 156,  29, 156,  28, 156,  27, 156,  26, 156,  25, 156,  24, 156,  23, 156,  22, 156,  21, 156,  20, 156,  19, 156,  18, 156,  17, 156,  16, 156,  15, 156,  14, 156,  13, 156,  12, 156,  11, 156,  10, 156,   9, 156,   8, 156,   7, 156,   6, 156,   5, 156,   4, 156,   3, 156,   2, 156,   1, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 156,   0, 143,  31, 143,  30, 143,  29, 143,  28, 143,  27, 143,  26, 143,  25, 143,  24, 143,  23, 143,  22, 143,  21, 143,  20, 143,  19, 143,  18, 143,  17, 143,  16, 143,  15, 143,  14, 143,  13, 143,  12, 143,  11, 143,  10, 143,   9, 143,   8, 143,   7, 143,   6, 143,   5, 143,   4, 143,   3, 143,   2, 143,   1, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 233,  31, 233,  30, 233,  29, 233,  28, 233,  27, 233,  26, 233,  25, 233,  24, 233,  23, 233,  22, 233,  21, 233,  20, 233,  19, 233,  18, 233,  17, 233,  16, 233,  15, 233,  14, 233,  13, 233,  12, 233,  11, 233,  10, 233,   9, 233,   8, 233,   7, 233,   6, 233,   5, 233,   4, 233,   3, 233,   2, 233,   1, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 233,   0, 200,  31, 200,  30, 200,  29, 200,  28, 200,  27, 200,  26, 200,  25, 200,  24, 200,  23, 200,  22, 200,  21, 200,  20, 200,  19, 200,  18, 200,  17, 200,  16, 200,  15,  91,  31,  91,  30,  91,  29,  91,  28,  91,  27,  91,  26,  91,  25,  91,  24,  91,  23,  91,  22,  91,  21,  91,  20,  91,  19,  91,  18,  91,  17,  91,  16,  35,  31,  35,  30,  35,  29,  35,  28,  35,  27,  35,  26,  35,  25,  35,  24,  70,  31,  70,  30,  70,  29,  70,  28,  70,  27,  70,  26,  70,  25,  70,  24,  70,  23,  70,  22,  70,  21,  70,  20,  70,  19,  70,  18,  70,  17,  70,  16,  70,  15,  70,  14,  70,  13,  70,  12,  70,  11,  70,  10,  70,   9,  70,   8,  70,   7,  70,   6,  70,   5,  70,   4,  70,   3,  70,   2,  70,   1,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0, 216,  31, 216,  30, 216,  29, 216,  28, 216,  27, 216,  26, 216,  25, 216,  24, 216,  23, 216,  22, 216,  21, 216,  20, 216,  19, 216,  18, 216,  17, 216,  16, 216,  15, 216,  14, 216,  13, 216,  12, 216,  11, 216,  10, 216,   9, 216,   8, 216,   7, 216,   6, 216,   5, 216,   4, 216,   3, 216,   2, 216,   1, 216,   0, 216,   0, 216,   0, 216,   0, 216,   0, 216,   0, 216,   0, 216,   0, 216,   0, 216,   0, 216,   0, 216,   0, 216,   0, 216,   0, 216,   0, 216,   0, 216,   0, 216,   0, 216,   0, 216,   0, 219,  31, 219,  30, 219,  29, 219,  28, 219,  27, 219,  26, 219,  25, 219,  24, 219,  23, 219,  22, 219,  21, 219,  20, 219,  19, 219,  18, 219,  17, 219,  16, 219,  15, 219,  14, 219,  13, 219,  12, 219,  11, 219,  10, 219,   9, 219,   8, 219,   7, 219,   6, 219,   5, 219,   4, 219,   3, 219,   2, 219,   1, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 219,   0, 176,  31, 176,  30, 176,  29, 176,  28, 176,  27, 176,  26, 176,  25, 176,  24, 176,  23, 176,  22, 176,  21, 176,  20, 176,  19, 176,  18, 176,  17, 176,  16, 176,  15, 176,  14, 176,  13, 176,  12, 176,  11, 176,  10, 176,   9, 176,   8, 176,   7, 176,   6, 176,   5, 176,   4, 176,   3, 176,   2, 176,   1, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 253,  31, 253,  30, 253,  29, 253,  28, 253,  27, 253,  26, 253,  25, 253,  24, 253,  23, 253,  22, 253,  21, 253,  20, 139,  31, 139,  30, 139,  29, 139,  28, 139,  27, 139,  26, 139,  25, 139,  24, 139,  23, 139,  22, 139,  21, 139,  20, 139,  19, 139,  18, 139,  17, 139,  16, 139,  15, 139,  14, 139,  13, 139,  12, 139,  11, 139,  10, 139,   9, 139,   8, 139,   7, 139,   6, 139,   5, 139,   4, 139,   3, 139,   2, 139,   1, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 139,   0, 170,  31, 170,  30, 170,  29, 170,  28, 170,  27, 170,  26, 170,  25, 170,  24, 170,  23, 170,  22, 170,  21, 191,  31, 191,  30, 191,  29, 191,  28, 191,  27, 191,  26, 191,  25, 191,  24, 191,  23, 191,  22, 191,  21, 191,  20, 191,  19, 191,  18, 191,  17, 191,  16, 191,  15, 191,  14, 191,  13, 191,  12, 191,  11, 191,  10, 191,   9, 191,   8, 191,   7, 191,   6, 191,   5, 191,   4, 191,   3, 191,   2, 191,   1, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 127,  31, 127,  30, 141,  31, 141,  30, 141,  29, 141,  28, 141,  27, 141,  26, 141,  25, 141,  24, 141,  23, 141,  22, 141,  21, 141,  20, 141,  19, 141,  18, 141,  17, 141,  16, 141,  15, 141,  14, 141,  13, 141,  12, 141,  11, 141,  10, 141,   9,  36,  31,  36,  30,  36,  29,  36,  28,  36,  27,  36,  26,  36,  25,  36,  24,  55,  31,  55,  30,  55,  29,  55,  28,  55,  27,  55,  26,  55,  25,  55,  24,  55,  23,  55,  22,  55,  21,  55,  20, 120,  31, 120,  30, 120,  29, 120,  28, 120,  27, 120,  26, 120,  25, 120,  24, 120,  23, 120,  22, 120,  21, 120,  20, 120,  19, 120,  18, 120,  17, 120,  16, 218,  31, 218,  30, 218,  29, 218,  28, 218,  27, 218,  26, 218,  25, 218,  24, 218,  23, 218,  22, 218,  21, 218,  20, 218,  19, 218,  18, 218,  17, 218,  16, 218,  15, 218,  14, 218,  13, 218,  12, 218,  11, 218,  10, 218,   9, 218,   8,  32,  31,  32,  30,  32,  29,  32,  28,  32,  27,  32,  26,  32,  25,  32,  24,  32,  23,  32,  22,  32,  21,  32,  20,  32,  19,  32,  18,  32,  17,  32,  16,  32,  15,  32,  14,  32,  13,  32,  12,  32,  11,  32,  10,  32,   9,  32,   8,  32,   7,  32,   6,  32,   5,  32,   4,  32,   3,  32,   2,  32,   1,  32,   0);
	constant SCENARIO_ADDRESS_25 : integer := 51246;


	--Scenario 26
	constant SCENARIO_LENGTH_26 : integer := 1006;
	type scenario_type_26 is array (0 to SCENARIO_LENGTH_26*2-1) of integer;
	signal scenario_input_26 : scenario_type_26 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  91,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 151,   0,   0,   0,  21,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  42,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 118,   0,   0,   0,   0,   0,  98,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  58,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 222,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 109,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 185,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  94,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  15,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 138,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 120,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 112,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  75,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  16,   0,   0,   0,   0,   0, 158,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  42,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 162,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  98,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  90,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 196,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 224,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  34,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  20,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 228,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_26  : scenario_type_26 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  91,  31,  91,  30,  91,  29,  91,  28,  91,  27,  91,  26,  91,  25,  91,  24,  91,  23,  91,  22,  91,  21,  91,  20,  91,  19,  91,  18,  91,  17,  91,  16,  91,  15, 151,  31, 151,  30,  21,  31,  21,  30,  21,  29,  21,  28,  21,  27,  21,  26,  21,  25,  21,  24,  21,  23,  21,  22,  21,  21,  21,  20,  21,  19,  21,  18,  21,  17,  21,  16,  21,  15,  21,  14,  21,  13,  21,  12,  21,  11,  21,  10,  21,   9,  21,   8,  21,   7,  21,   6,  21,   5,  21,   4,  21,   3,  21,   2,  21,   1,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  21,   0,  42,  31,  42,  30,  42,  29,  42,  28,  42,  27,  42,  26,  42,  25,  42,  24,  42,  23,  42,  22,  42,  21,  42,  20,  42,  19,  42,  18,  42,  17,  42,  16,  42,  15,  42,  14,  42,  13,  42,  12, 118,  31, 118,  30, 118,  29,  98,  31,  98,  30,  98,  29,  98,  28,  98,  27,  98,  26,  98,  25,  98,  24,  98,  23,  98,  22,  58,  31,  58,  30,  58,  29,  58,  28,  58,  27,  58,  26,  58,  25,  58,  24,  58,  23,  58,  22,  58,  21,  58,  20,  58,  19,  58,  18,  58,  17,  58,  16,  58,  15,  58,  14,  58,  13,  58,  12,  58,  11,  58,  10,  58,   9,  58,   8,  58,   7,  58,   6,  58,   5,  58,   4,  58,   3,  58,   2,  58,   1,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0,  58,   0, 222,  31, 222,  30, 222,  29, 222,  28, 222,  27, 222,  26, 222,  25, 222,  24, 222,  23, 222,  22, 222,  21, 222,  20, 222,  19, 222,  18, 222,  17, 222,  16, 222,  15, 222,  14, 222,  13, 222,  12, 222,  11, 222,  10, 222,   9, 222,   8, 222,   7, 222,   6, 222,   5, 222,   4, 222,   3, 222,   2, 222,   1, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 222,   0, 109,  31, 109,  30, 109,  29, 109,  28, 109,  27, 109,  26, 109,  25, 109,  24, 109,  23, 109,  22, 109,  21, 109,  20, 109,  19, 109,  18, 109,  17, 109,  16, 109,  15, 109,  14, 109,  13, 109,  12, 109,  11, 109,  10, 109,   9, 109,   8, 109,   7, 109,   6, 109,   5, 109,   4, 109,   3, 109,   2, 185,  31, 185,  30, 185,  29, 185,  28, 185,  27, 185,  26, 185,  25, 185,  24, 185,  23, 185,  22, 185,  21, 185,  20, 185,  19, 185,  18, 185,  17, 185,  16,  94,  31,  94,  30,  94,  29,  94,  28,  94,  27,  94,  26,  94,  25,  94,  24,  94,  23,  94,  22,  94,  21,  94,  20,  94,  19,  15,  31,  15,  30,  15,  29,  15,  28,  15,  27,  15,  26,  15,  25,  15,  24,  15,  23,  15,  22,  15,  21,  15,  20,  15,  19,  15,  18,  15,  17,  15,  16,  15,  15,  15,  14,  15,  13,  15,  12,  15,  11,  15,  10,  15,   9,  15,   8,  15,   7,  15,   6,  15,   5,  15,   4,  15,   3,  15,   2,  15,   1,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0, 138,  31, 138,  30, 138,  29, 138,  28, 138,  27, 138,  26, 138,  25, 138,  24, 138,  23, 138,  22, 138,  21, 138,  20, 138,  19, 138,  18, 138,  17, 120,  31, 120,  30, 120,  29, 120,  28, 120,  27, 120,  26, 120,  25, 120,  24, 120,  23, 120,  22, 120,  21, 120,  20, 120,  19, 120,  18, 120,  17, 120,  16, 120,  15, 120,  14, 120,  13, 120,  12, 120,  11, 120,  10, 120,   9, 120,   8, 120,   7, 120,   6, 120,   5, 120,   4, 120,   3, 120,   2, 120,   1, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 112,  31, 112,  30, 112,  29, 112,  28, 112,  27, 112,  26, 112,  25, 112,  24, 112,  23,  75,  31,  75,  30,  75,  29,  75,  28,  75,  27,  75,  26,  75,  25,  75,  24,  75,  23,  75,  22,  75,  21,  75,  20,  75,  19,  75,  18,  75,  17,  75,  16,  75,  15,  75,  14,  75,  13,  75,  12,  75,  11,  75,  10,  75,   9,  75,   8,  75,   7,  75,   6,  75,   5,  75,   4,  75,   3,  75,   2,  75,   1,  75,   0,  75,   0,  75,   0,  75,   0,  75,   0,  75,   0,  75,   0,  75,   0,  75,   0,  75,   0,  75,   0,  75,   0,  75,   0,  75,   0,  75,   0,  75,   0,  75,   0,  75,   0,  75,   0,  75,   0,  75,   0,  75,   0,  16,  31,  16,  30,  16,  29, 158,  31, 158,  30, 158,  29, 158,  28, 158,  27, 158,  26, 158,  25, 158,  24, 158,  23, 158,  22, 158,  21, 158,  20, 158,  19, 158,  18, 158,  17, 158,  16, 158,  15, 158,  14, 158,  13, 158,  12, 158,  11, 158,  10, 158,   9, 158,   8, 158,   7, 158,   6, 158,   5, 158,   4, 158,   3, 158,   2, 158,   1, 158,   0, 158,   0, 158,   0, 158,   0, 158,   0, 158,   0, 158,   0, 158,   0,  42,  31,  42,  30,  42,  29,  42,  28,  42,  27,  42,  26,  42,  25, 162,  31, 162,  30, 162,  29, 162,  28, 162,  27, 162,  26, 162,  25, 162,  24, 162,  23, 162,  22, 162,  21, 162,  20, 162,  19, 162,  18, 162,  17, 162,  16, 162,  15, 162,  14, 162,  13, 162,  12, 162,  11, 162,  10, 162,   9, 162,   8, 162,   7, 162,   6, 162,   5, 162,   4, 162,   3, 162,   2, 162,   1, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0,  98,  31,  98,  30,  98,  29,  98,  28,  98,  27,  98,  26,  98,  25,  98,  24,  98,  23,  98,  22,  98,  21,  98,  20,  98,  19,  98,  18,  98,  17,  98,  16,  98,  15,  98,  14,  98,  13,  98,  12,  98,  11,  98,  10,  98,   9,  90,  31,  90,  30,  90,  29,  90,  28,  90,  27,  90,  26,  90,  25,  90,  24,  90,  23,  90,  22,  90,  21,  90,  20,  90,  19,  90,  18,  90,  17,  90,  16,  90,  15,  90,  14,  90,  13,  90,  12,  90,  11, 196,  31, 196,  30, 196,  29, 196,  28, 196,  27, 196,  26, 196,  25, 196,  24, 196,  23, 196,  22, 196,  21, 196,  20, 196,  19, 196,  18, 196,  17, 196,  16, 196,  15, 196,  14, 224,  31, 224,  30, 224,  29, 224,  28, 224,  27, 224,  26, 224,  25, 224,  24, 224,  23, 224,  22, 224,  21, 224,  20, 224,  19, 224,  18, 224,  17, 224,  16, 224,  15, 224,  14, 224,  13, 224,  12, 224,  11, 224,  10, 224,   9, 224,   8, 224,   7, 224,   6, 224,   5, 224,   4, 224,   3, 224,   2, 224,   1, 224,   0, 224,   0, 224,   0, 224,   0, 224,   0, 224,   0, 224,   0, 224,   0, 224,   0, 224,   0, 224,   0, 224,   0, 224,   0, 224,   0, 224,   0, 224,   0,  34,  31,  34,  30,  34,  29,  34,  28,  34,  27,  34,  26,  34,  25,  34,  24,  34,  23,  34,  22,  34,  21,  34,  20,  34,  19,  34,  18,  34,  17,  34,  16,  34,  15,  34,  14,  34,  13,  34,  12,  34,  11,  34,  10,  34,   9,  34,   8,  34,   7,  34,   6,  34,   5,  34,   4,  34,   3,  34,   2,  34,   1,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0,  20,  31,  20,  30,  20,  29,  20,  28,  20,  27,  20,  26,  20,  25,  20,  24,  20,  23,  20,  22,  20,  21,  20,  20,  20,  19,  20,  18,  20,  17,  20,  16,  20,  15,  20,  14,  20,  13,  20,  12,  20,  11,  20,  10,  20,   9,  20,   8,  20,   7,  20,   6,  20,   5,  20,   4,  20,   3,  20,   2,  20,   1,  20,   0,  20,   0,  20,   0,  20,   0,  20,   0,  20,   0,  20,   0,  20,   0,  20,   0,  20,   0,  20,   0,  20,   0,  20,   0,  20,   0,  20,   0,  20,   0,  20,   0,  20,   0,  20,   0,  20,   0, 228,  31, 228,  30, 228,  29, 228,  28, 228,  27, 228,  26, 228,  25, 228,  24, 228,  23, 228,  22, 228,  21);
	constant SCENARIO_ADDRESS_26 : integer := 53269;


	--Scenario 27
	constant SCENARIO_LENGTH_27 : integer := 985;
	type scenario_type_27 is array (0 to SCENARIO_LENGTH_27*2-1) of integer;
	signal scenario_input_27 : scenario_type_27 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 199,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 146,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  10,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 176,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  60,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 140,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   2,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 176,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   6,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   2,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 120,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  13,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  73,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 180,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 242,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  91,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 104,   0,   0,   0,   0,   0,   0,   0,   0,   0, 117,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  95,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 146,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  39,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  51,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 245,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 131,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 239,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 213,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  97,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 200,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  91,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  31,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_27  : scenario_type_27 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 199,  31, 199,  30, 199,  29, 199,  28, 199,  27, 199,  26, 199,  25, 199,  24, 199,  23, 199,  22, 199,  21, 199,  20, 199,  19, 199,  18, 199,  17, 199,  16, 199,  15, 199,  14, 199,  13, 199,  12, 199,  11, 199,  10, 199,   9, 199,   8, 199,   7, 199,   6, 199,   5, 199,   4, 199,   3, 199,   2, 199,   1, 199,   0, 199,   0, 199,   0, 199,   0, 199,   0, 199,   0, 199,   0, 199,   0, 199,   0, 199,   0, 199,   0, 199,   0, 199,   0, 199,   0, 199,   0, 199,   0, 199,   0, 146,  31, 146,  30, 146,  29, 146,  28, 146,  27, 146,  26, 146,  25, 146,  24, 146,  23, 146,  22, 146,  21, 146,  20, 146,  19, 146,  18, 146,  17, 146,  16, 146,  15, 146,  14, 146,  13, 146,  12,  10,  31,  10,  30,  10,  29,  10,  28,  10,  27,  10,  26,  10,  25,  10,  24,  10,  23,  10,  22,  10,  21,  10,  20,  10,  19,  10,  18,  10,  17,  10,  16,  10,  15,  10,  14,  10,  13,  10,  12,  10,  11,  10,  10,  10,   9,  10,   8,  10,   7,  10,   6,  10,   5,  10,   4,  10,   3,  10,   2,  10,   1,  10,   0, 176,  31, 176,  30, 176,  29, 176,  28, 176,  27, 176,  26, 176,  25, 176,  24, 176,  23, 176,  22, 176,  21, 176,  20, 176,  19, 176,  18, 176,  17, 176,  16, 176,  15, 176,  14, 176,  13, 176,  12, 176,  11, 176,  10, 176,   9, 176,   8, 176,   7, 176,   6, 176,   5, 176,   4, 176,   3, 176,   2, 176,   1, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0, 176,   0,  60,  31,  60,  30,  60,  29,  60,  28,  60,  27,  60,  26,  60,  25,  60,  24,  60,  23,  60,  22,  60,  21,  60,  20,  60,  19,  60,  18,  60,  17,  60,  16,  60,  15,  60,  14,  60,  13,  60,  12,  60,  11,  60,  10,  60,   9,  60,   8,  60,   7,  60,   6,  60,   5,  60,   4,  60,   3,  60,   2,  60,   1,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0,  60,   0, 140,  31, 140,  30, 140,  29, 140,  28, 140,  27, 140,  26, 140,  25, 140,  24, 140,  23, 140,  22, 140,  21, 140,  20, 140,  19, 140,  18, 140,  17, 140,  16, 140,  15, 140,  14, 140,  13, 140,  12, 140,  11, 140,  10, 140,   9, 140,   8, 140,   7, 140,   6, 140,   5, 140,   4, 140,   3, 140,   2, 140,   1, 140,   0, 140,   0, 140,   0, 140,   0, 140,   0, 140,   0, 140,   0, 140,   0, 140,   0, 140,   0, 140,   0, 140,   0, 140,   0, 140,   0, 140,   0, 140,   0, 140,   0,   2,  31,   2,  30,   2,  29,   2,  28,   2,  27,   2,  26,   2,  25,   2,  24,   2,  23,   2,  22,   2,  21,   2,  20,   2,  19,   2,  18,   2,  17,   2,  16,   2,  15,   2,  14,   2,  13,   2,  12,   2,  11,   2,  10,   2,   9,   2,   8,   2,   7,   2,   6,   2,   5,   2,   4,   2,   3,   2,   2, 176,  31, 176,  30, 176,  29, 176,  28, 176,  27, 176,  26, 176,  25, 176,  24, 176,  23, 176,  22, 176,  21, 176,  20, 176,  19, 176,  18, 176,  17,   6,  31,   6,  30,   6,  29,   6,  28,   6,  27,   6,  26,   6,  25,   6,  24,   6,  23,   6,  22,   6,  21,   6,  20,   6,  19,   6,  18,   6,  17,   6,  16,   6,  15,   6,  14,   6,  13,   2,  31,   2,  30,   2,  29,   2,  28,   2,  27,   2,  26,   2,  25,   2,  24,   2,  23,   2,  22,   2,  21,   2,  20,   2,  19,   2,  18,   2,  17,   2,  16,   2,  15,   2,  14,   2,  13,   2,  12,   2,  11,   2,  10,   2,   9,   2,   8,   2,   7,   2,   6,   2,   5,   2,   4,   2,   3,   2,   2,   2,   1, 120,  31, 120,  30, 120,  29, 120,  28, 120,  27, 120,  26, 120,  25, 120,  24, 120,  23, 120,  22, 120,  21, 120,  20, 120,  19, 120,  18, 120,  17, 120,  16, 120,  15, 120,  14, 120,  13, 120,  12, 120,  11, 120,  10, 120,   9, 120,   8, 120,   7, 120,   6, 120,   5, 120,   4, 120,   3, 120,   2, 120,   1, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0, 120,   0,  13,  31,  13,  30,  13,  29,  13,  28,  13,  27,  13,  26,  13,  25,  13,  24,  13,  23,  13,  22,  13,  21,  73,  31,  73,  30,  73,  29,  73,  28,  73,  27,  73,  26,  73,  25,  73,  24,  73,  23,  73,  22,  73,  21,  73,  20,  73,  19,  73,  18,  73,  17,  73,  16,  73,  15,  73,  14,  73,  13,  73,  12,  73,  11,  73,  10,  73,   9,  73,   8,  73,   7, 180,  31, 180,  30, 180,  29, 180,  28, 180,  27, 180,  26, 180,  25, 180,  24, 180,  23, 180,  22, 180,  21, 180,  20, 180,  19, 180,  18, 180,  17, 180,  16, 180,  15, 180,  14, 180,  13, 180,  12, 180,  11, 180,  10, 180,   9, 180,   8, 180,   7, 180,   6, 180,   5, 180,   4, 180,   3, 180,   2, 180,   1, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 242,  31, 242,  30, 242,  29, 242,  28, 242,  27, 242,  26, 242,  25, 242,  24, 242,  23, 242,  22, 242,  21, 242,  20, 242,  19, 242,  18, 242,  17, 242,  16, 242,  15, 242,  14, 242,  13, 242,  12, 242,  11, 242,  10, 242,   9, 242,   8, 242,   7, 242,   6, 242,   5, 242,   4, 242,   3, 242,   2, 242,   1, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0, 242,   0,  91,  31,  91,  30,  91,  29,  91,  28,  91,  27,  91,  26,  91,  25,  91,  24,  91,  23,  91,  22,  91,  21,  91,  20,  91,  19,  91,  18,  91,  17,  91,  16,  91,  15,  91,  14,  91,  13,  91,  12,  91,  11,  91,  10,  91,   9,  91,   8,  91,   7,  91,   6,  91,   5,  91,   4, 104,  31, 104,  30, 104,  29, 104,  28, 104,  27, 117,  31, 117,  30, 117,  29, 117,  28, 117,  27, 117,  26, 117,  25, 117,  24, 117,  23, 117,  22, 117,  21,  95,  31,  95,  30,  95,  29,  95,  28,  95,  27,  95,  26,  95,  25,  95,  24,  95,  23,  95,  22, 146,  31, 146,  30, 146,  29, 146,  28, 146,  27, 146,  26, 146,  25, 146,  24, 146,  23, 146,  22, 146,  21, 146,  20, 146,  19, 146,  18, 146,  17, 146,  16, 146,  15, 146,  14, 146,  13, 146,  12, 146,  11, 146,  10, 146,   9, 146,   8, 146,   7, 146,   6, 146,   5, 146,   4, 146,   3, 146,   2, 146,   1, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0, 146,   0,  39,  31,  39,  30,  39,  29,  39,  28,  39,  27,  39,  26,  39,  25,  39,  24,  39,  23,  39,  22,  39,  21,  39,  20,  39,  19,  39,  18,  39,  17,  39,  16,  39,  15,  39,  14,  39,  13,  39,  12,  39,  11,  39,  10,  39,   9,  39,   8,  39,   7,  51,  31,  51,  30,  51,  29,  51,  28,  51,  27,  51,  26,  51,  25,  51,  24,  51,  23,  51,  22,  51,  21,  51,  20,  51,  19,  51,  18,  51,  17,  51,  16,  51,  15,  51,  14,  51,  13,  51,  12,  51,  11,  51,  10,  51,   9,  51,   8,  51,   7,  51,   6,  51,   5,  51,   4,  51,   3,  51,   2,  51,   1, 245,  31, 245,  30, 245,  29, 245,  28, 245,  27, 245,  26, 245,  25, 245,  24, 245,  23, 245,  22, 245,  21, 245,  20, 245,  19, 245,  18, 245,  17, 245,  16, 245,  15, 245,  14, 245,  13, 245,  12, 245,  11, 245,  10, 245,   9, 245,   8, 245,   7, 245,   6, 245,   5, 245,   4, 245,   3, 245,   2, 245,   1, 245,   0, 245,   0, 245,   0, 245,   0, 245,   0, 131,  31, 131,  30, 131,  29, 131,  28, 131,  27, 131,  26, 131,  25, 131,  24, 131,  23, 131,  22, 131,  21, 131,  20, 131,  19, 131,  18, 131,  17, 131,  16, 131,  15, 131,  14, 131,  13, 239,  31, 239,  30, 239,  29, 239,  28, 239,  27, 239,  26, 239,  25, 239,  24, 239,  23, 239,  22, 239,  21, 239,  20, 239,  19, 239,  18, 239,  17, 239,  16, 239,  15, 239,  14, 239,  13, 239,  12, 239,  11, 239,  10, 239,   9, 239,   8, 239,   7, 239,   6, 239,   5, 239,   4, 239,   3, 239,   2, 239,   1, 239,   0, 239,   0, 239,   0, 239,   0, 213,  31, 213,  30, 213,  29, 213,  28, 213,  27, 213,  26, 213,  25, 213,  24,  97,  31,  97,  30,  97,  29,  97,  28,  97,  27,  97,  26,  97,  25,  97,  24,  97,  23,  97,  22,  97,  21,  97,  20, 200,  31, 200,  30, 200,  29, 200,  28, 200,  27, 200,  26, 200,  25, 200,  24, 200,  23, 200,  22, 200,  21, 200,  20, 200,  19, 200,  18, 200,  17, 200,  16, 200,  15, 200,  14, 200,  13, 200,  12, 200,  11, 200,  10, 200,   9, 200,   8, 200,   7, 200,   6, 200,   5, 200,   4, 200,   3, 200,   2, 200,   1, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0,  91,  31,  91,  30,  91,  29,  91,  28,  91,  27,  91,  26,  91,  25,  91,  24,  91,  23,  91,  22,  91,  21,  91,  20,  91,  19,  91,  18,  91,  17,  91,  16,  91,  15,  91,  14,  91,  13,  91,  12,  91,  11,  91,  10,  91,   9,  91,   8,  91,   7,  91,   6,  91,   5,  91,   4,  91,   3,  91,   2,  91,   1,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  91,   0,  31,  31,  31,  30,  31,  29,  31,  28,  31,  27,  31,  26);
	constant SCENARIO_ADDRESS_27 : integer := 55353;


	--Scenario 28
	constant SCENARIO_LENGTH_28 : integer := 984;
	type scenario_type_28 is array (0 to SCENARIO_LENGTH_28*2-1) of integer;
	signal scenario_input_28 : scenario_type_28 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 203,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 118,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  29,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 206,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 170,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 147,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 197,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 190,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 181,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 229,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 199,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 191,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  64,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 243,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 127,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 247,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 187,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 129,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 255,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 180,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 129,   0, 133,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 197,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  19,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  74,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 217,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 217,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 251,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 200,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_28  : scenario_type_28 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 203,  31, 203,  30, 203,  29, 203,  28, 203,  27, 203,  26, 203,  25, 203,  24, 203,  23, 203,  22, 203,  21, 203,  20, 203,  19, 203,  18, 203,  17, 203,  16, 203,  15, 203,  14, 203,  13, 203,  12, 203,  11, 203,  10, 203,   9, 203,   8, 203,   7, 203,   6, 203,   5, 203,   4, 203,   3, 203,   2, 203,   1, 203,   0, 203,   0, 203,   0, 203,   0, 203,   0, 203,   0, 203,   0, 203,   0, 203,   0, 203,   0, 203,   0, 203,   0, 203,   0, 118,  31, 118,  30, 118,  29, 118,  28, 118,  27, 118,  26, 118,  25, 118,  24, 118,  23, 118,  22, 118,  21, 118,  20, 118,  19, 118,  18, 118,  17, 118,  16, 118,  15, 118,  14, 118,  13, 118,  12, 118,  11, 118,  10, 118,   9, 118,   8, 118,   7, 118,   6, 118,   5, 118,   4, 118,   3, 118,   2, 118,   1, 118,   0,  29,  31,  29,  30,  29,  29,  29,  28,  29,  27,  29,  26,  29,  25,  29,  24,  29,  23,  29,  22,  29,  21,  29,  20,  29,  19,  29,  18,  29,  17,  29,  16,  29,  15,  29,  14,  29,  13,  29,  12,  29,  11, 206,  31, 206,  30, 206,  29, 206,  28, 206,  27, 206,  26, 206,  25, 206,  24, 206,  23, 206,  22, 206,  21, 206,  20, 206,  19, 206,  18, 206,  17, 206,  16, 206,  15, 206,  14, 206,  13, 206,  12, 206,  11, 206,  10, 206,   9, 206,   8, 206,   7, 206,   6, 206,   5, 206,   4, 206,   3, 206,   2, 206,   1, 206,   0, 206,   0, 206,   0, 206,   0, 206,   0, 206,   0, 206,   0, 206,   0, 206,   0, 206,   0, 206,   0, 206,   0, 206,   0, 206,   0, 206,   0, 206,   0, 206,   0, 206,   0, 170,  31, 170,  30, 170,  29, 170,  28, 170,  27, 170,  26, 170,  25, 170,  24, 170,  23, 170,  22, 170,  21, 170,  20, 170,  19, 170,  18, 170,  17, 170,  16, 170,  15, 170,  14, 170,  13, 170,  12, 170,  11, 170,  10, 170,   9, 170,   8, 170,   7, 170,   6, 170,   5, 170,   4, 170,   3, 170,   2, 170,   1, 170,   0, 170,   0, 170,   0, 170,   0, 170,   0, 170,   0, 170,   0, 170,   0, 170,   0, 170,   0, 170,   0, 170,   0, 170,   0, 170,   0, 170,   0, 170,   0, 170,   0, 170,   0, 170,   0, 170,   0, 170,   0, 147,  31, 147,  30, 147,  29, 147,  28, 147,  27, 147,  26, 147,  25, 147,  24, 147,  23, 197,  31, 197,  30, 197,  29, 197,  28, 197,  27, 197,  26, 190,  31, 190,  30, 190,  29, 190,  28, 190,  27, 190,  26, 190,  25, 190,  24, 190,  23, 190,  22, 190,  21, 190,  20, 190,  19, 190,  18, 190,  17, 190,  16, 190,  15, 190,  14, 190,  13, 190,  12, 190,  11, 190,  10, 190,   9, 190,   8, 190,   7, 190,   6, 190,   5, 190,   4, 190,   3, 190,   2, 190,   1, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 190,   0, 181,  31, 181,  30, 181,  29, 181,  28, 181,  27, 181,  26, 181,  25, 181,  24, 181,  23, 181,  22, 181,  21, 181,  20, 181,  19, 181,  18, 181,  17, 181,  16, 181,  15, 181,  14, 229,  31, 229,  30, 229,  29, 229,  28, 229,  27, 229,  26, 229,  25, 229,  24, 229,  23, 229,  22, 229,  21, 229,  20, 229,  19, 229,  18, 229,  17, 229,  16, 229,  15, 229,  14, 229,  13, 229,  12, 229,  11, 229,  10, 229,   9, 229,   8, 229,   7, 229,   6, 229,   5, 229,   4, 229,   3, 229,   2, 199,  31, 199,  30, 199,  29, 199,  28, 199,  27, 199,  26, 199,  25, 199,  24, 199,  23, 199,  22, 191,  31, 191,  30, 191,  29, 191,  28, 191,  27, 191,  26, 191,  25, 191,  24, 191,  23, 191,  22, 191,  21, 191,  20, 191,  19, 191,  18, 191,  17, 191,  16, 191,  15, 191,  14, 191,  13, 191,  12, 191,  11, 191,  10, 191,   9, 191,   8, 191,   7, 191,   6, 191,   5, 191,   4, 191,   3, 191,   2, 191,   1, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0, 191,   0,  64,  31,  64,  30,  64,  29,  64,  28,  64,  27,  64,  26,  64,  25,  64,  24,  64,  23,  64,  22,  64,  21,  64,  20,  64,  19,  64,  18,  64,  17,  64,  16,  64,  15,  64,  14,  64,  13,  64,  12,  64,  11,  64,  10,  64,   9,  64,   8,  64,   7,  64,   6,  64,   5,  64,   4,  64,   3,  64,   2,  64,   1,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0, 243,  31, 243,  30, 243,  29, 243,  28, 243,  27, 243,  26, 243,  25, 243,  24, 243,  23, 243,  22, 243,  21, 243,  20, 243,  19, 243,  18, 243,  17, 243,  16, 243,  15, 243,  14, 243,  13, 243,  12, 243,  11, 243,  10, 243,   9, 243,   8, 243,   7, 243,   6, 243,   5, 243,   4, 243,   3, 243,   2, 243,   1, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 243,   0, 127,  31, 127,  30, 127,  29, 127,  28, 127,  27, 127,  26, 127,  25, 127,  24, 127,  23, 127,  22, 127,  21, 127,  20, 127,  19, 127,  18, 127,  17, 127,  16, 127,  15, 127,  14, 127,  13, 127,  12, 127,  11, 127,  10, 127,   9, 127,   8, 127,   7, 127,   6, 127,   5, 127,   4, 127,   3, 127,   2, 127,   1, 247,  31, 247,  30, 247,  29, 247,  28, 247,  27, 247,  26, 247,  25, 247,  24, 247,  23, 247,  22, 247,  21, 247,  20, 247,  19, 247,  18, 247,  17, 247,  16, 247,  15, 247,  14, 247,  13, 247,  12, 247,  11, 247,  10, 247,   9, 247,   8, 247,   7, 247,   6, 247,   5, 247,   4, 247,   3, 247,   2, 247,   1, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 187,  31, 187,  30, 187,  29, 187,  28, 187,  27, 187,  26, 187,  25, 187,  24, 187,  23, 187,  22, 187,  21, 187,  20, 187,  19, 187,  18, 129,  31, 129,  30, 129,  29, 129,  28, 129,  27, 129,  26, 129,  25, 129,  24, 129,  23, 129,  22, 129,  21, 129,  20, 129,  19, 129,  18, 129,  17, 129,  16, 129,  15, 129,  14, 129,  13, 129,  12, 129,  11, 129,  10, 129,   9, 129,   8, 129,   7, 129,   6, 129,   5, 129,   4, 129,   3, 129,   2, 129,   1, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 129,   0, 255,  31, 255,  30, 255,  29, 255,  28, 255,  27, 255,  26, 255,  25, 255,  24, 255,  23, 255,  22, 255,  21, 255,  20, 255,  19, 255,  18, 255,  17, 255,  16, 255,  15, 255,  14, 255,  13, 255,  12, 255,  11, 255,  10, 255,   9, 255,   8, 255,   7, 255,   6, 255,   5, 255,   4, 255,   3, 255,   2, 255,   1, 255,   0, 255,   0, 255,   0, 180,  31, 180,  30, 180,  29, 180,  28, 180,  27, 180,  26, 180,  25, 180,  24, 180,  23, 180,  22, 180,  21, 180,  20, 180,  19, 180,  18, 180,  17, 180,  16, 180,  15, 180,  14, 180,  13, 180,  12, 180,  11, 180,  10, 180,   9, 180,   8, 180,   7, 180,   6, 180,   5, 180,   4, 180,   3, 180,   2, 180,   1, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 180,   0, 129,  31, 133,  31, 133,  30, 133,  29, 133,  28, 133,  27, 133,  26, 133,  25, 133,  24, 133,  23, 133,  22, 133,  21, 133,  20, 133,  19, 197,  31, 197,  30, 197,  29, 197,  28, 197,  27, 197,  26, 197,  25, 197,  24, 197,  23, 197,  22, 197,  21, 197,  20, 197,  19, 197,  18, 197,  17, 197,  16, 197,  15, 197,  14, 197,  13, 197,  12, 197,  11, 197,  10, 197,   9, 197,   8, 197,   7, 197,   6, 197,   5, 197,   4, 197,   3, 197,   2, 197,   1, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0, 197,   0,  19,  31,  19,  30,  19,  29,  19,  28,  19,  27,  19,  26,  19,  25,  19,  24,  19,  23,  19,  22,  19,  21,  19,  20,  19,  19,  19,  18,  19,  17,  19,  16,  19,  15,  19,  14,  19,  13,  19,  12,  19,  11,  19,  10,  19,   9,  19,   8,  19,   7,  19,   6,  19,   5,  19,   4,  19,   3,  19,   2,  19,   1,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  19,   0,  74,  31,  74,  30,  74,  29,  74,  28,  74,  27,  74,  26,  74,  25,  74,  24,  74,  23,  74,  22,  74,  21,  74,  20,  74,  19,  74,  18,  74,  17,  74,  16,  74,  15,  74,  14,  74,  13,  74,  12,  74,  11,  74,  10,  74,   9,  74,   8,  74,   7,  74,   6,  74,   5,  74,   4,  74,   3,  74,   2,  74,   1,  74,   0,  74,   0,  74,   0,  74,   0,  74,   0,  74,   0,  74,   0,  74,   0,  74,   0,  74,   0,  74,   0,  74,   0,  74,   0,  74,   0,  74,   0,  74,   0,  74,   0,  74,   0, 217,  31, 217,  30, 217,  29, 217,  28, 217,  27, 217,  26, 217,  25, 217,  24, 217,  23, 217,  22, 217,  21, 217,  20, 217,  19, 217,  18, 217,  17, 217,  16, 217,  15, 217,  14, 217,  13, 217,  12, 217,  11, 217,  10, 217,   9, 217,   8, 217,   7, 217,   6, 217,   5, 217,   4, 217,  31, 217,  30, 217,  29, 217,  28, 217,  27, 217,  26, 217,  25, 217,  24, 217,  23, 217,  22, 217,  21, 217,  20, 217,  19, 217,  18, 217,  17, 217,  16, 217,  15, 251,  31, 251,  30, 251,  29, 251,  28, 251,  27, 251,  26, 251,  25, 251,  24, 251,  23, 251,  22, 251,  21, 251,  20, 251,  19, 251,  18, 251,  17, 251,  16, 251,  15, 251,  14, 200,  31, 200,  30, 200,  29, 200,  28, 200,  27, 200,  26, 200,  25, 200,  24, 200,  23, 200,  22, 200,  21, 200,  20, 200,  19, 200,  18, 200,  17, 200,  16, 200,  15, 200,  14, 200,  13, 200,  12, 200,  11, 200,  10, 200,   9, 200,   8, 200,   7, 200,   6, 200,   5, 200,   4, 200,   3, 200,   2, 200,   1, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0, 200,   0);
	constant SCENARIO_ADDRESS_28 : integer := 57400;


	--Scenario 29
	constant SCENARIO_LENGTH_29 : integer := 1016;
	type scenario_type_29 is array (0 to SCENARIO_LENGTH_29*2-1) of integer;
	signal scenario_input_29 : scenario_type_29 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 235,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  50,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  27,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 253,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 143,   0,   0,   0,   0,   0,   0,   0, 123,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 107,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 143,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  46,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  29,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  17,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  99,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 182,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 194,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 125,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 162,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  79,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  74,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 125,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  96,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 183,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 168,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 201,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  25,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 190,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 132,   0,   0,   0,   0,   0,   0,   0,   0,   0, 156,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 139,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_29  : scenario_type_29 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 235,  31, 235,  30, 235,  29, 235,  28, 235,  27, 235,  26, 235,  25, 235,  24, 235,  23, 235,  22, 235,  21, 235,  20, 235,  19, 235,  18, 235,  17, 235,  16, 235,  15, 235,  14, 235,  13, 235,  12, 235,  11, 235,  10, 235,   9, 235,   8, 235,   7, 235,   6, 235,   5, 235,   4, 235,   3, 235,   2, 235,   1, 235,   0, 235,   0, 235,   0, 235,   0, 235,   0, 235,   0, 235,   0, 235,   0, 235,   0, 235,   0, 235,   0, 235,   0, 235,   0, 235,   0, 235,   0, 235,   0, 235,   0, 235,   0,  50,  31,  50,  30,  50,  29,  50,  28,  50,  27,  50,  26,  50,  25,  50,  24,  50,  23,  50,  22,  50,  21,  50,  20,  50,  19,  50,  18,  50,  17,  50,  16,  50,  15,  50,  14,  50,  13,  50,  12,  50,  11,  50,  10,  50,   9,  50,   8,  50,   7,  50,   6,  50,   5,  50,   4,  50,   3,  50,   2,  50,   1,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  50,   0,  27,  31,  27,  30,  27,  29,  27,  28,  27,  27,  27,  26,  27,  25,  27,  24,  27,  23,  27,  22,  27,  21,  27,  20, 253,  31, 253,  30, 253,  29, 253,  28, 253,  27, 253,  26, 253,  25, 253,  24, 253,  23, 253,  22, 253,  21, 253,  20, 253,  19, 253,  18, 253,  17, 253,  16, 253,  15, 253,  14, 253,  13, 253,  12, 253,  11, 253,  10, 253,   9, 253,   8, 253,   7, 253,   6, 253,   5, 253,   4, 253,   3, 253,   2, 253,   1, 253,   0, 253,   0, 253,   0, 253,   0, 253,   0, 253,   0, 253,   0, 253,   0, 253,   0, 143,  31, 143,  30, 143,  29, 143,  28, 123,  31, 123,  30, 123,  29, 123,  28, 123,  27, 123,  26, 123,  25, 123,  24, 123,  23, 123,  22, 123,  21, 123,  20, 123,  19, 123,  18, 123,  17, 123,  16, 123,  15, 123,  14, 123,  13, 123,  12, 123,  11, 123,  10, 123,   9, 123,   8, 123,   7, 123,   6, 123,   5, 123,   4, 123,   3, 123,   2, 123,   1, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 123,   0, 107,  31, 107,  30, 107,  29, 107,  28, 107,  27, 107,  26, 107,  25, 107,  24, 107,  23, 107,  22, 107,  21, 107,  20, 107,  19, 107,  18, 107,  17, 107,  16, 107,  15, 107,  14, 107,  13, 107,  12, 107,  11, 107,  10, 107,   9, 107,   8, 107,   7, 107,   6, 107,   5, 107,   4, 107,   3, 107,   2, 107,   1, 107,   0, 107,   0, 107,   0, 107,   0, 107,   0, 107,   0, 107,   0, 107,   0, 107,   0, 107,   0, 107,   0, 107,   0, 107,   0, 107,   0, 143,  31, 143,  30, 143,  29, 143,  28, 143,  27, 143,  26, 143,  25, 143,  24, 143,  23, 143,  22, 143,  21, 143,  20, 143,  19, 143,  18, 143,  17, 143,  16, 143,  15, 143,  14, 143,  13, 143,  12, 143,  11, 143,  10, 143,   9, 143,   8, 143,   7, 143,   6, 143,   5, 143,   4, 143,   3, 143,   2, 143,   1, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0, 143,   0,  46,  31,  46,  30,  46,  29,  46,  28,  46,  27,  46,  26,  46,  25,  46,  24,  46,  23,  46,  22,  46,  21,  46,  20,  46,  19,  46,  18,  46,  17,  46,  16,  46,  15,  46,  14,  46,  13,  46,  12,  46,  11,  46,  10,  46,   9,  46,   8,  46,   7,  46,   6,  46,   5,  46,   4,  46,   3,  46,   2,  46,   1,  46,   0,  46,   0,  46,   0,  29,  31,  29,  30,  29,  29,  29,  28,  29,  27,  29,  26,  29,  25,  29,  24,  29,  23,  29,  22,  29,  21,  29,  20,  29,  19,  29,  18,  29,  17,  29,  16,  29,  15,  29,  14,  29,  13,  29,  12,  29,  11,  29,  10,  29,   9,  29,   8,  29,   7,  29,   6,  29,   5,  29,   4,  29,   3,  29,   2,  29,   1,  29,   0,  29,   0,  29,   0,  29,   0,  29,   0,  29,   0,  29,   0,  29,   0,  29,   0,  29,   0,  29,   0,  29,   0,  29,   0,  17,  31,  17,  30,  17,  29,  17,  28,  17,  27,  17,  26,  17,  25,  17,  24,  17,  23,  17,  22,  17,  21,  17,  20,  17,  19,  17,  18,  17,  17,  17,  16,  17,  15,  17,  14,  17,  13,  17,  12,  17,  11,  17,  10,  17,   9,  17,   8,  17,   7,  17,   6,  17,   5,  17,   4,  17,   3,  17,   2,  17,   1,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  17,   0,  99,  31,  99,  30,  99,  29,  99,  28,  99,  27,  99,  26,  99,  25,  99,  24,  99,  23,  99,  22,  99,  21,  99,  20,  99,  19,  99,  18,  99,  17,  99,  16,  99,  15,  99,  14,  99,  13,  99,  12,  99,  11,  99,  10,  99,   9,  99,   8,  99,   7,  99,   6,  99,   5,  99,   4,  99,   3,  99,   2,  99,   1,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0, 182,  31, 182,  30, 182,  29, 182,  28, 182,  27, 182,  26, 182,  25, 182,  24, 182,  23, 182,  22, 182,  21, 182,  20, 182,  19, 182,  18, 182,  17, 182,  16, 182,  15, 182,  14, 182,  13, 182,  12, 182,  11, 182,  10, 182,   9, 194,  31, 194,  30, 194,  29, 194,  28, 194,  27, 194,  26, 194,  25, 194,  24, 194,  23, 194,  22, 194,  21, 194,  20, 194,  19, 194,  18, 194,  17, 194,  16, 194,  15, 194,  14, 194,  13, 194,  12, 194,  11, 194,  10, 194,   9, 194,   8, 194,   7, 194,   6, 194,   5, 194,   4, 194,   3, 194,   2, 194,   1, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 194,   0, 125,  31, 125,  30, 125,  29, 125,  28, 125,  27, 125,  26, 125,  25, 125,  24, 125,  23, 125,  22, 125,  21, 125,  20, 125,  19, 125,  18, 125,  17, 125,  16, 125,  15, 125,  14, 125,  13, 125,  12, 125,  11, 125,  10, 125,   9, 125,   8, 125,   7, 125,   6, 125,   5, 125,   4, 125,   3, 125,   2, 125,   1, 125,   0, 125,   0, 125,   0, 125,   0, 162,  31, 162,  30, 162,  29, 162,  28, 162,  27, 162,  26, 162,  25, 162,  24, 162,  23, 162,  22, 162,  21, 162,  20, 162,  19, 162,  18, 162,  17, 162,  16, 162,  15, 162,  14, 162,  13, 162,  12, 162,  11, 162,  10, 162,   9, 162,   8, 162,   7, 162,   6, 162,   5, 162,   4, 162,   3, 162,   2, 162,   1, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0, 162,   0,  79,  31,  79,  30,  79,  29,  79,  28,  79,  27,  79,  26,  79,  25,  79,  24,  79,  23,  79,  22,  74,  31,  74,  30,  74,  29,  74,  28,  74,  27,  74,  26,  74,  25,  74,  24,  74,  23,  74,  22,  74,  21,  74,  20,  74,  19,  74,  18,  74,  17,  74,  16,  74,  15,  74,  14,  74,  13,  74,  12,  74,  11,  74,  10,  74,   9,  74,   8,  74,   7,  74,   6,  74,   5,  74,   4,  74,   3,  74,   2,  74,   1,  74,   0,  74,   0,  74,   0, 125,  31, 125,  30, 125,  29, 125,  28, 125,  27, 125,  26, 125,  25, 125,  24, 125,  23, 125,  22, 125,  21, 125,  20, 125,  19, 125,  18, 125,  17, 125,  16, 125,  15, 125,  14, 125,  13, 125,  12, 125,  11, 125,  10, 125,   9, 125,   8, 125,   7, 125,   6, 125,   5, 125,   4, 125,   3, 125,   2, 125,   1, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0, 125,   0,  96,  31,  96,  30,  96,  29,  96,  28,  96,  27,  96,  26,  96,  25,  96,  24,  96,  23,  96,  22,  96,  21,  96,  20,  96,  19,  96,  18,  96,  17,  96,  16,  96,  15,  96,  14,  96,  13,  96,  12,  96,  11,  96,  10,  96,   9,  96,   8,  96,   7,  96,   6,  96,   5,  96,   4, 183,  31, 183,  30, 183,  29, 183,  28, 183,  27, 183,  26, 183,  25, 183,  24, 183,  23, 183,  22, 183,  21, 183,  20, 183,  19, 183,  18, 183,  17, 183,  16, 183,  15, 183,  14, 183,  13, 183,  12, 183,  11, 183,  10, 183,   9, 183,   8, 183,   7, 183,   6, 183,   5, 183,   4, 168,  31, 168,  30, 168,  29, 168,  28, 168,  27, 168,  26, 168,  25, 168,  24, 168,  23, 168,  22, 168,  21, 168,  20, 168,  19, 168,  18, 168,  17, 168,  16, 168,  15, 168,  14, 168,  13, 168,  12, 168,  11, 168,  10, 168,   9, 168,   8, 168,   7, 168,   6, 168,   5, 168,   4, 201,  31, 201,  30, 201,  29, 201,  28, 201,  27, 201,  26, 201,  25, 201,  24,  25,  31,  25,  30,  25,  29,  25,  28,  25,  27,  25,  26,  25,  25,  25,  24,  25,  23,  25,  22,  25,  21,  25,  20,  25,  19,  25,  18,  25,  17,  25,  16,  25,  15,  25,  14,  25,  13,  25,  12,  25,  11,  25,  10,  25,   9,  25,   8,  25,   7,  25,   6,  25,   5,  25,   4,  25,   3,  25,   2,  25,   1,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0,  25,   0, 190,  31, 190,  30, 190,  29, 190,  28, 190,  27, 190,  26, 190,  25, 190,  24, 190,  23, 190,  22, 190,  21, 190,  20, 190,  19, 190,  18, 190,  17, 190,  16, 190,  15, 190,  14, 190,  13, 190,  12, 190,  11, 190,  10, 190,   9, 190,   8, 190,   7, 190,   6, 190,   5, 190,   4, 190,   3, 190,   2, 190,   1, 132,  31, 132,  30, 132,  29, 132,  28, 132,  27, 156,  31, 156,  30, 156,  29, 156,  28, 156,  27, 156,  26, 156,  25, 156,  24, 156,  23, 156,  22, 156,  21, 139,  31, 139,  30, 139,  29, 139,  28, 139,  27, 139,  26, 139,  25, 139,  24, 139,  23, 139,  22, 139,  21, 139,  20);
	constant SCENARIO_ADDRESS_29 : integer := 59396;


	--Scenario 30
	constant SCENARIO_LENGTH_30 : integer := 1005;
	type scenario_type_30 is array (0 to SCENARIO_LENGTH_30*2-1) of integer;
	signal scenario_input_30 : scenario_type_30 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  14,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  70,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  18,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 105,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 119,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  70,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 170,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 220,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  43,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 160,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 202,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  46,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 227,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  32,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  64,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 110,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  88,   0,   0,   0,   0,   0, 142,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 131,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  39,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  34,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 185,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 173,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 145,   0,   0,   0,  32,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  16,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  55,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  60,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_30  : scenario_type_30 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  14,  31,  14,  30,  14,  29,  14,  28,  14,  27,  14,  26,  14,  25,  14,  24,  14,  23,  14,  22,  14,  21,  14,  20,  14,  19,  14,  18,  14,  17,  14,  16,  14,  15,  14,  14,  14,  13,  14,  12,  14,  11,  14,  10,  14,   9,  14,   8,  14,   7,  14,   6,  14,   5,  14,   4,  14,   3,  14,   2,  14,   1,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  14,   0,  70,  31,  70,  30,  70,  29,  70,  28,  70,  27,  70,  26,  70,  25,  70,  24,  70,  23,  70,  22,  70,  21,  70,  20,  70,  19,  70,  18,  70,  17,  70,  16,  70,  15,  70,  14,  70,  13,  70,  12,  70,  11,  70,  10,  70,   9,  70,   8,  70,   7,  70,   6,  70,   5,  70,   4,  70,   3,  70,   2,  70,   1,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0,  18,  31,  18,  30,  18,  29,  18,  28,  18,  27,  18,  26,  18,  25,  18,  24,  18,  23,  18,  22,  18,  21,  18,  20,  18,  19,  18,  18,  18,  17,  18,  16,  18,  15,  18,  14,  18,  13,  18,  12,  18,  11,  18,  10,  18,   9,  18,   8,  18,   7,  18,   6,  18,   5,  18,   4,  18,   3,  18,   2,  18,   1,  18,   0,  18,   0,  18,   0,  18,   0,  18,   0,  18,   0,  18,   0,  18,   0,  18,   0, 105,  31, 105,  30, 105,  29, 105,  28, 105,  27, 105,  26, 105,  25, 105,  24, 105,  23, 105,  22, 105,  21, 105,  20, 105,  19, 105,  18, 105,  17, 105,  16, 105,  15, 105,  14, 105,  13, 105,  12, 105,  11, 105,  10, 105,   9, 105,   8, 105,   7, 105,   6, 105,   5, 105,   4, 105,   3, 105,   2, 105,   1, 105,   0, 105,   0, 105,   0, 105,   0, 105,   0, 105,   0, 105,   0, 105,   0, 105,   0, 105,   0, 105,   0, 105,   0, 105,   0, 105,   0, 105,   0, 119,  31, 119,  30, 119,  29, 119,  28, 119,  27, 119,  26, 119,  25, 119,  24, 119,  23, 119,  22, 119,  21, 119,  20, 119,  19, 119,  18, 119,  17, 119,  16, 119,  15, 119,  14, 119,  13, 119,  12, 119,  11, 119,  10, 119,   9, 119,   8, 119,   7, 119,   6, 119,   5, 119,   4, 119,   3, 119,   2, 119,   1, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0, 119,   0,  70,  31,  70,  30,  70,  29,  70,  28,  70,  27,  70,  26,  70,  25,  70,  24,  70,  23,  70,  22,  70,  21,  70,  20,  70,  19,  70,  18,  70,  17,  70,  16,  70,  15,  70,  14,  70,  13,  70,  12,  70,  11,  70,  10,  70,   9,  70,   8,  70,   7,  70,   6,  70,   5,  70,   4,  70,   3,  70,   2,  70,   1,  70,   0,  70,   0,  70,   0,  70,   0,  70,   0, 170,  31, 170,  30, 170,  29, 170,  28, 170,  27, 170,  26, 170,  25, 170,  24, 170,  23, 170,  22, 170,  21, 170,  20, 170,  19, 170,  18, 170,  17, 170,  16, 170,  15, 170,  14, 170,  13, 170,  12, 170,  11, 170,  10, 220,  31, 220,  30, 220,  29, 220,  28, 220,  27, 220,  26, 220,  25, 220,  24, 220,  23, 220,  22, 220,  21, 220,  20, 220,  19, 220,  18, 220,  17, 220,  16, 220,  15, 220,  14, 220,  13, 220,  12, 220,  11, 220,  10, 220,   9, 220,   8, 220,   7, 220,   6, 220,   5, 220,   4, 220,   3, 220,   2, 220,   1, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0, 220,   0,  43,  31,  43,  30,  43,  29,  43,  28,  43,  27,  43,  26,  43,  25,  43,  24,  43,  23,  43,  22,  43,  21,  43,  20,  43,  19,  43,  18,  43,  17,  43,  16,  43,  15,  43,  14, 160,  31, 160,  30, 160,  29, 160,  28, 160,  27, 160,  26, 160,  25, 160,  24, 160,  23, 160,  22, 160,  21, 160,  20, 160,  19, 160,  18, 160,  17, 160,  16, 160,  15, 160,  14, 160,  13, 160,  12, 202,  31, 202,  30, 202,  29, 202,  28, 202,  27, 202,  26, 202,  25, 202,  24, 202,  23, 202,  22, 202,  21, 202,  20, 202,  19, 202,  18, 202,  17, 202,  16, 202,  15, 202,  14, 202,  13, 202,  12, 202,  11, 202,  10, 202,   9, 202,   8, 202,   7, 202,   6, 202,   5, 202,   4, 202,   3, 202,   2, 202,   1, 202,   0, 202,   0, 202,   0, 202,   0, 202,   0, 202,   0, 202,   0, 202,   0, 202,   0, 202,   0,  46,  31,  46,  30,  46,  29,  46,  28,  46,  27,  46,  26,  46,  25,  46,  24,  46,  23,  46,  22,  46,  21,  46,  20,  46,  19,  46,  18,  46,  17,  46,  16,  46,  15,  46,  14,  46,  13,  46,  12,  46,  11,  46,  10,  46,   9,  46,   8,  46,   7,  46,   6,  46,   5,  46,   4,  46,   3,  46,   2,  46,   1,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0,  46,   0, 227,  31, 227,  30, 227,  29, 227,  28, 227,  27, 227,  26, 227,  25, 227,  24, 227,  23, 227,  22, 227,  21, 227,  20, 227,  19, 227,  18, 227,  17, 227,  16, 227,  15, 227,  14, 227,  13, 227,  12, 227,  11,  32,  31,  32,  30,  32,  29,  32,  28,  32,  27,  32,  26,  32,  25,  32,  24,  32,  23,  32,  22,  32,  21,  32,  20,  32,  19,  32,  18,  32,  17,  32,  16,  32,  15,  32,  14,  32,  13,  32,  12,  32,  11,  32,  10,  32,   9,  32,   8,  32,   7,  32,   6,  32,   5,  32,   4,  32,   3,  32,   2,  32,   1,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  32,   0,  64,  31,  64,  30,  64,  29,  64,  28,  64,  27,  64,  26,  64,  25,  64,  24,  64,  23,  64,  22,  64,  21,  64,  20,  64,  19,  64,  18,  64,  17,  64,  16,  64,  15,  64,  14,  64,  13,  64,  12,  64,  11,  64,  10,  64,   9,  64,   8,  64,   7,  64,   6,  64,   5,  64,   4,  64,   3,  64,   2,  64,   1,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0,  64,   0, 110,  31, 110,  30, 110,  29, 110,  28, 110,  27, 110,  26, 110,  25, 110,  24, 110,  23, 110,  22, 110,  21, 110,  20, 110,  19, 110,  18, 110,  17, 110,  16, 110,  15, 110,  14, 110,  13, 110,  12, 110,  11, 110,  10, 110,   9, 110,   8, 110,   7, 110,   6, 110,   5, 110,   4, 110,   3, 110,   2, 110,   1, 110,   0, 110,   0, 110,   0, 110,   0, 110,   0, 110,   0, 110,   0,  88,  31,  88,  30,  88,  29, 142,  31, 142,  30, 142,  29, 142,  28, 142,  27, 142,  26, 142,  25, 142,  24, 142,  23, 142,  22, 142,  21, 142,  20, 142,  19, 142,  18, 142,  17, 142,  16, 142,  15, 142,  14, 142,  13, 142,  12, 142,  11, 142,  10, 142,   9, 142,   8, 142,   7, 142,   6, 142,   5, 142,   4, 142,   3, 142,   2, 142,   1, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 142,   0, 131,  31, 131,  30, 131,  29, 131,  28, 131,  27, 131,  26, 131,  25, 131,  24, 131,  23, 131,  22, 131,  21, 131,  20, 131,  19, 131,  18, 131,  17, 131,  16, 131,  15, 131,  14, 131,  13, 131,  12, 131,  11, 131,  10,  39,  31,  39,  30,  39,  29,  39,  28,  39,  27,  39,  26,  39,  25,  39,  24,  39,  23,  39,  22,  39,  21,  39,  20,  39,  19,  39,  18,  39,  17,  39,  16,  39,  15,  34,  31,  34,  30,  34,  29,  34,  28,  34,  27,  34,  26,  34,  25,  34,  24,  34,  23,  34,  22,  34,  21,  34,  20,  34,  19,  34,  18,  34,  17,  34,  16,  34,  15,  34,  14,  34,  13,  34,  12,  34,  11,  34,  10,  34,   9,  34,   8,  34,   7,  34,   6,  34,   5,  34,   4,  34,   3,  34,   2,  34,   1,  34,   0,  34,   0,  34,   0,  34,   0,  34,   0, 185,  31, 185,  30, 185,  29, 185,  28, 185,  27, 185,  26, 185,  25, 185,  24, 185,  23, 185,  22, 185,  21, 185,  20, 185,  19, 185,  18, 185,  17, 185,  16, 185,  15, 185,  14, 185,  13, 185,  12, 185,  11, 185,  10, 185,   9, 185,   8, 185,   7, 185,   6, 185,   5, 185,   4, 185,   3, 185,   2, 185,   1, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 185,   0, 173,  31, 173,  30, 173,  29, 173,  28, 173,  27, 173,  26, 173,  25, 173,  24, 173,  23, 173,  22, 173,  21, 173,  20, 173,  19, 173,  18, 173,  17, 173,  16, 173,  15, 173,  14, 173,  13, 173,  12, 173,  11, 173,  10, 173,   9, 173,   8, 173,   7, 173,   6, 173,   5, 173,   4, 173,   3, 173,   2, 173,   1, 173,   0, 173,   0, 145,  31, 145,  30,  32,  31,  32,  30,  32,  29,  32,  28,  32,  27,  32,  26,  16,  31,  16,  30,  16,  29,  16,  28,  16,  27,  16,  26,  16,  25,  16,  24,  16,  23,  16,  22,  16,  21,  16,  20,  16,  19,  16,  18,  16,  17,  16,  16,  16,  15,  16,  14,  16,  13,  16,  12,  16,  11,  16,  10,  16,   9,  16,   8,  16,   7,  16,   6,  16,   5,  16,   4,  16,   3,  16,   2,  16,   1,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  16,   0,  55,  31,  55,  30,  55,  29,  55,  28,  55,  27,  55,  26,  55,  25,  55,  24,  55,  23,  55,  22,  55,  21,  55,  20,  55,  19,  55,  18,  55,  17,  55,  16,  55,  15,  55,  14,  55,  13,  55,  12,  55,  11,  55,  10,  55,   9,  60,  31,  60,  30,  60,  29,  60,  28,  60,  27,  60,  26,  60,  25,  60,  24,  60,  23);
	constant SCENARIO_ADDRESS_30 : integer := 61472;


	--Scenario 31
	constant SCENARIO_LENGTH_31 : integer := 986;
	type scenario_type_31 is array (0 to SCENARIO_LENGTH_31*2-1) of integer;
	signal scenario_input_31 : scenario_type_31 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 233,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 164,   0,   0,   0, 216,   0,   0,   0,   0,   0,  69,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  40,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  67,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 188,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  22,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   7,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 254,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 232,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 202,   0,   0,   0,   0,   0,  42,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 249,   0,   0,   0,   0,   0, 227,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  90,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  15,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 144,   0,   0,   0,   0,   0,   0,   0, 129,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 247,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 183,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 250,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  32,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  95,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  99,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 133,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 229,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,  67,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 180,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 141,   0,   0,   0, 118,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 171,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0);
	signal scenario_full_31  : scenario_type_31 := (0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0,   0, 233,  31, 233,  30, 233,  29, 233,  28, 233,  27, 233,  26, 233,  25, 233,  24, 233,  23, 233,  22, 233,  21, 233,  20, 233,  19, 233,  18, 233,  17, 233,  16, 233,  15, 233,  14, 233,  13, 164,  31, 164,  30, 216,  31, 216,  30, 216,  29,  69,  31,  69,  30,  69,  29,  69,  28,  69,  27,  69,  26,  69,  25,  69,  24,  69,  23,  69,  22,  69,  21,  69,  20,  69,  19,  40,  31,  40,  30,  40,  29,  40,  28,  40,  27,  40,  26,  40,  25,  40,  24,  40,  23,  40,  22,  40,  21,  40,  20,  40,  19,  40,  18,  40,  17,  40,  16,  40,  15,  40,  14,  40,  13,  40,  12,  40,  11,  40,  10,  40,   9,  40,   8,  40,   7,  40,   6,  40,   5,  40,   4,  40,   3,  40,   2,  40,   1,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  40,   0,  67,  31,  67,  30,  67,  29,  67,  28,  67,  27,  67,  26,  67,  25,  67,  24,  67,  23,  67,  22,  67,  21,  67,  20,  67,  19,  67,  18,  67,  17,  67,  16,  67,  15,  67,  14,  67,  13,  67,  12,  67,  11,  67,  10,  67,   9,  67,   8,  67,   7,  67,   6,  67,   5,  67,   4,  67,   3,  67,   2,  67,   1,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0, 188,  31, 188,  30, 188,  29, 188,  28, 188,  27, 188,  26, 188,  25, 188,  24, 188,  23, 188,  22, 188,  21, 188,  20, 188,  19, 188,  18, 188,  17, 188,  16, 188,  15, 188,  14, 188,  13, 188,  12, 188,  11, 188,  10, 188,   9, 188,   8, 188,   7, 188,   6, 188,   5, 188,   4, 188,   3, 188,   2, 188,   1, 188,   0, 188,   0,  22,  31,  22,  30,  22,  29,  22,  28,  22,  27,  22,  26,  22,  25,  22,  24,  22,  23,  22,  22,  22,  21,  22,  20,  22,  19,  22,  18,  22,  17,  22,  16,  22,  15,  22,  14,  22,  13,  22,  12,  22,  11,  22,  10,  22,   9,  22,   8,  22,   7,  22,   6,  22,   5,  22,   4,  22,   3,  22,   2,  22,   1,   7,  31,   7,  30,   7,  29,   7,  28,   7,  27,   7,  26,   7,  25,   7,  24,   7,  23,   7,  22,   7,  21,   7,  20,   7,  19,   7,  18,   7,  17,   7,  16,   7,  15,   7,  14,   7,  13,   7,  12,   7,  11,   7,  10,   7,   9,   7,   8,   7,   7,   7,   6,   7,   5,   7,   4, 254,  31, 254,  30, 254,  29, 254,  28, 254,  27, 254,  26, 254,  25, 254,  24, 254,  23, 254,  22, 232,  31, 232,  30, 232,  29, 232,  28, 232,  27, 232,  26, 232,  25, 232,  24, 232,  23, 232,  22, 232,  21, 232,  20, 232,  19, 232,  18, 232,  17, 232,  16, 202,  31, 202,  30, 202,  29,  42,  31,  42,  30,  42,  29,  42,  28,  42,  27,  42,  26,  42,  25,  42,  24,  42,  23,  42,  22,  42,  21,  42,  20,  42,  19,  42,  18,  42,  17,  42,  16,  42,  15,  42,  14,  42,  13,  42,  12,  42,  11,  42,  10,  42,   9,  42,   8,  42,   7,  42,   6,  42,   5, 249,  31, 249,  30, 249,  29, 227,  31, 227,  30, 227,  29, 227,  28, 227,  27, 227,  26, 227,  25, 227,  24, 227,  23, 227,  22, 227,  21, 227,  20, 227,  19, 227,  18, 227,  17,  90,  31,  90,  30,  90,  29,  90,  28,  90,  27,  90,  26,  90,  25,  90,  24,  90,  23,  90,  22,  90,  21,  90,  20,  90,  19,  90,  18,  90,  17,  90,  16,  90,  15,  90,  14,  90,  13,  90,  12,  90,  11,  90,  10,  90,   9,  90,   8,  90,   7,  90,   6,  90,   5,  90,   4,  90,   3,  90,   2,  15,  31,  15,  30,  15,  29,  15,  28,  15,  27,  15,  26,  15,  25,  15,  24,  15,  23,  15,  22,  15,  21,  15,  20,  15,  19,  15,  18,  15,  17,  15,  16,  15,  15,  15,  14,  15,  13,  15,  12,  15,  11,  15,  10,  15,   9,  15,   8,  15,   7,  15,   6,  15,   5,  15,   4,  15,   3,  15,   2,  15,   1,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0,  15,   0, 144,  31, 144,  30, 144,  29, 144,  28, 129,  31, 129,  30, 129,  29, 129,  28, 129,  27, 129,  26, 129,  25, 129,  24, 129,  23, 129,  22, 129,  21, 129,  20, 129,  19, 129,  18, 247,  31, 247,  30, 247,  29, 247,  28, 247,  27, 247,  26, 247,  25, 247,  24, 247,  23, 247,  22, 247,  21, 247,  20, 247,  19, 247,  18, 247,  17, 247,  16, 247,  15, 247,  14, 247,  13, 247,  12, 247,  11, 247,  10, 247,   9, 247,   8, 247,   7, 247,   6, 247,   5, 247,   4, 247,   3, 247,   2, 247,   1, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 247,   0, 183,  31, 183,  30, 183,  29, 183,  28, 183,  27, 183,  26, 183,  25, 183,  24, 183,  23, 183,  22, 183,  21, 183,  20, 183,  19, 183,  18, 183,  17, 183,  16, 183,  15, 183,  14, 183,  13, 183,  12, 183,  11, 183,  10, 183,   9, 183,   8, 183,   7, 183,   6, 183,   5, 183,   4, 183,   3, 183,   2, 183,   1, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 183,   0, 250,  31, 250,  30, 250,  29, 250,  28, 250,  27, 250,  26, 250,  25, 250,  24, 250,  23, 250,  22, 250,  21, 250,  20, 250,  19, 250,  18, 250,  17, 250,  16, 250,  15, 250,  14, 250,  13, 250,  12, 250,  11, 250,  10, 250,   9, 250,   8, 250,   7, 250,   6, 250,   5, 250,   4, 250,   3, 250,   2, 250,   1, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0, 250,   0,  32,  31,  32,  30,  32,  29,  32,  28,  32,  27,  32,  26,  32,  25,  32,  24,  32,  23,  32,  22,  32,  21,  32,  20,  32,  19,  32,  18,  32,  17,  32,  16,  32,  15,  32,  14,  32,  13,  32,  12,  32,  11,  32,  10,  32,   9,  32,   8,  32,   7,  32,   6,  32,   5,  32,   4,  32,   3,  32,   2,  32,   1,  32,   0,  95,  31,  95,  30,  95,  29,  95,  28,  95,  27,  95,  26,  95,  25,  95,  24,  95,  23,  95,  22,  95,  21,  95,  20,  95,  19,  95,  18,  95,  17,  95,  16,  95,  15,  95,  14,  95,  13,  95,  12,  95,  11,  95,  10,  95,   9,  95,   8,  95,   7,  95,   6,  95,   5,  95,   4,  95,   3,  95,   2,  95,   1,  95,   0,  95,   0,  99,  31,  99,  30,  99,  29,  99,  28,  99,  27,  99,  26,  99,  25,  99,  24,  99,  23,  99,  22,  99,  21,  99,  20,  99,  19,  99,  18,  99,  17,  99,  16,  99,  15,  99,  14,  99,  13,  99,  12,  99,  11,  99,  10,  99,   9,  99,   8,  99,   7,  99,   6,  99,   5,  99,   4,  99,   3,  99,   2,  99,   1,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0,  99,   0, 133,  31, 133,  30, 133,  29, 133,  28, 133,  27, 133,  26, 133,  25, 133,  24, 133,  23, 133,  22, 133,  21, 133,  20, 133,  19, 133,  18, 133,  17, 133,  16, 133,  15, 133,  14, 133,  13, 133,  12, 133,  11, 133,  10, 133,   9, 133,   8, 133,   7, 133,   6, 133,   5, 133,   4, 133,   3, 229,  31, 229,  30, 229,  29, 229,  28, 229,  27, 229,  26, 229,  25, 229,  24, 229,  23, 229,  22, 229,  21, 229,  20, 229,  19, 229,  18, 229,  17, 229,  16, 229,  15, 229,  14, 229,  13, 229,  12, 229,  11, 229,  10, 229,   9, 229,   8, 229,   7, 229,   6, 229,   5, 229,   4, 229,   3, 229,   2, 229,   1, 229,   0, 229,   0, 229,   0, 229,   0, 229,   0, 229,   0, 229,   0,  67,  31,  67,  30,  67,  29,  67,  28,  67,  27,  67,  26,  67,  25,  67,  24,  67,  23,  67,  22,  67,  21,  67,  20,  67,  19,  67,  18,  67,  17,  67,  16,  67,  15,  67,  14,  67,  13,  67,  12,  67,  11,  67,  10,  67,   9,  67,   8,  67,   7,  67,   6,  67,   5,  67,   4,  67,   3,  67,   2,  67,   1,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0,  67,   0, 180,  31, 180,  30, 180,  29, 180,  28, 180,  27, 180,  26, 180,  25, 180,  24, 180,  23, 180,  22, 180,  21, 180,  20, 180,  19, 180,  18, 141,  31, 141,  30, 118,  31, 118,  30, 118,  29, 118,  28, 118,  27, 118,  26, 118,  25, 118,  24, 118,  23, 118,  22, 118,  21, 118,  20, 118,  19, 118,  18, 118,  17, 118,  16, 118,  15, 118,  14, 118,  13, 118,  12, 118,  11, 118,  10, 118,   9, 118,   8, 118,   7, 118,   6, 118,   5, 118,   4, 118,   3, 118,   2, 118,   1, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 118,   0, 171,  31, 171,  30, 171,  29, 171,  28, 171,  27, 171,  26, 171,  25, 171,  24, 171,  23, 171,  22, 171,  21, 171,  20, 171,  19, 171,  18, 171,  17, 171,  16, 171,  15, 171,  14, 171,  13, 171,  12, 171,  11, 171,  10, 171,   9, 171,   8, 171,   7, 171,   6, 171,   5, 171,   4, 171,   3, 171,   2, 171,   1, 171,   0);
	constant SCENARIO_ADDRESS_31 : integer := 63534;

-- End Scenario Definition

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory 

-- Memory Initialization

		--Scenario 0
		for i in 0 to SCENARIO_LENGTH_0*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_0+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_0(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 1
		for i in 0 to SCENARIO_LENGTH_1*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_1+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_1(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 2
		for i in 0 to SCENARIO_LENGTH_2*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_2+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_2(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 3
		for i in 0 to SCENARIO_LENGTH_3*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_3+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_3(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 4
		for i in 0 to SCENARIO_LENGTH_4*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_4+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_4(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 5
		for i in 0 to SCENARIO_LENGTH_5*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_5+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_5(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 6
		for i in 0 to SCENARIO_LENGTH_6*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_6+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_6(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 7
		for i in 0 to SCENARIO_LENGTH_7*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_7+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_7(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 8
		for i in 0 to SCENARIO_LENGTH_8*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_8+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_8(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 9
		for i in 0 to SCENARIO_LENGTH_9*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_9+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_9(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 10
		for i in 0 to SCENARIO_LENGTH_10*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_10+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_10(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 11
		for i in 0 to SCENARIO_LENGTH_11*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_11+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_11(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 12
		for i in 0 to SCENARIO_LENGTH_12*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_12+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_12(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 13
		for i in 0 to SCENARIO_LENGTH_13*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_13+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_13(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 14
		for i in 0 to SCENARIO_LENGTH_14*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_14+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_14(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 15
		for i in 0 to SCENARIO_LENGTH_15*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_15+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_15(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 16
		for i in 0 to SCENARIO_LENGTH_16*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_16+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_16(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 17
		for i in 0 to SCENARIO_LENGTH_17*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_17+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_17(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 18
		for i in 0 to SCENARIO_LENGTH_18*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_18+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_18(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 19
		for i in 0 to SCENARIO_LENGTH_19*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_19+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_19(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 20
		for i in 0 to SCENARIO_LENGTH_20*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_20+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_20(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 21
		for i in 0 to SCENARIO_LENGTH_21*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_21+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_21(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 22
		for i in 0 to SCENARIO_LENGTH_22*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_22+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_22(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 23
		for i in 0 to SCENARIO_LENGTH_23*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_23+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_23(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 24
		for i in 0 to SCENARIO_LENGTH_24*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_24+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_24(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 25
		for i in 0 to SCENARIO_LENGTH_25*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_25+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_25(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 26
		for i in 0 to SCENARIO_LENGTH_26*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_26+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_26(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 27
		for i in 0 to SCENARIO_LENGTH_27*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_27+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_27(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 28
		for i in 0 to SCENARIO_LENGTH_28*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_28+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_28(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 29
		for i in 0 to SCENARIO_LENGTH_29*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_29+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_29(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 30
		for i in 0 to SCENARIO_LENGTH_30*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_30+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_30(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;


		--Scenario 31
		for i in 0 to SCENARIO_LENGTH_31*2-1 loop
			init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_31+i, 16));
			init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_31(i),8));
			init_o_mem_en  <= '1';
			init_o_mem_we  <= '1';
			wait until rising_edge(tb_clk); 
		end loop;

-- End Memory Initialization
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

-- Computation

	--Scenario 0
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_0, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_0, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 1
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_1, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_1, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 2
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_2, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_2, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 3
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_3, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_3, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 4
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_4, 16));
	tb_k   <= std_logic_vector(to_unsigned(0, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 5
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_5, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_5, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 6
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_6, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_6, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 7
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_7, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_7, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 8
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_8, 16));
	tb_k   <= std_logic_vector(to_unsigned(0, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 9
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_9, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_9, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 10
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_10, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_10, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 11
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_11, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_11, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 12
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_12, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_12, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 13
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_13, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_13, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 14
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_14, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_14, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 15
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_15, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_15, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 16
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_16, 16));
	tb_k   <= std_logic_vector(to_unsigned(0, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 17
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_17, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_17, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 18
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_18, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_18, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 19
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_19, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_19, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 20
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_20, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_20, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 21
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_21, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_21, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 22
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_22, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_22, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 23
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_23, 16));
	tb_k   <= std_logic_vector(to_unsigned(0, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 24
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_24, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_24, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 25
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_25, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_25, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 26
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_26, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_26, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 27
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_27, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_27, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 28
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_28, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_28, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 29
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_29, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_29, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 30
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_30, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_30, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);

	--Scenario 31
	tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_31, 16));
	tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_31, 10));

	tb_start <= '1';

	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	wait for 5 ns;

	tb_start <= '0';
	wait until falling_edge(tb_done);
-- End Computation
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
		
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;

-- Test

	--Scenario 0
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_0*2-1 loop
	assert RAM(SCENARIO_ADDRESS_0+i) = std_logic_vector(to_unsigned(scenario_full_0(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_0(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_0+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 1
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_1*2-1 loop
	assert RAM(SCENARIO_ADDRESS_1+i) = std_logic_vector(to_unsigned(scenario_full_1(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_1(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_1+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 2
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_2*2-1 loop
	assert RAM(SCENARIO_ADDRESS_2+i) = std_logic_vector(to_unsigned(scenario_full_2(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_2(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_2+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 3
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_3*2-1 loop
	assert RAM(SCENARIO_ADDRESS_3+i) = std_logic_vector(to_unsigned(scenario_full_3(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_3(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_3+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 4
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_4*2-1 loop
	assert RAM(SCENARIO_ADDRESS_4+i) = std_logic_vector(to_unsigned(scenario_full_4(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_4(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_4+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 5
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_5*2-1 loop
	assert RAM(SCENARIO_ADDRESS_5+i) = std_logic_vector(to_unsigned(scenario_full_5(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_5(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_5+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 6
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_6*2-1 loop
	assert RAM(SCENARIO_ADDRESS_6+i) = std_logic_vector(to_unsigned(scenario_full_6(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_6(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_6+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 7
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_7*2-1 loop
	assert RAM(SCENARIO_ADDRESS_7+i) = std_logic_vector(to_unsigned(scenario_full_7(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_7(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_7+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 8
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_8*2-1 loop
	assert RAM(SCENARIO_ADDRESS_8+i) = std_logic_vector(to_unsigned(scenario_full_8(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_8(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_8+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 9
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_9*2-1 loop
	assert RAM(SCENARIO_ADDRESS_9+i) = std_logic_vector(to_unsigned(scenario_full_9(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_9(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_9+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 10
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_10*2-1 loop
	assert RAM(SCENARIO_ADDRESS_10+i) = std_logic_vector(to_unsigned(scenario_full_10(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_10(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_10+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 11
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_11*2-1 loop
	assert RAM(SCENARIO_ADDRESS_11+i) = std_logic_vector(to_unsigned(scenario_full_11(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_11(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_11+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 12
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_12*2-1 loop
	assert RAM(SCENARIO_ADDRESS_12+i) = std_logic_vector(to_unsigned(scenario_full_12(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_12(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_12+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 13
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_13*2-1 loop
	assert RAM(SCENARIO_ADDRESS_13+i) = std_logic_vector(to_unsigned(scenario_full_13(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_13(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_13+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 14
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_14*2-1 loop
	assert RAM(SCENARIO_ADDRESS_14+i) = std_logic_vector(to_unsigned(scenario_full_14(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_14(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_14+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 15
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_15*2-1 loop
	assert RAM(SCENARIO_ADDRESS_15+i) = std_logic_vector(to_unsigned(scenario_full_15(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_15(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_15+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 16
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_16*2-1 loop
	assert RAM(SCENARIO_ADDRESS_16+i) = std_logic_vector(to_unsigned(scenario_full_16(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_16(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_16+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 17
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_17*2-1 loop
	assert RAM(SCENARIO_ADDRESS_17+i) = std_logic_vector(to_unsigned(scenario_full_17(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_17(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_17+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 18
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_18*2-1 loop
	assert RAM(SCENARIO_ADDRESS_18+i) = std_logic_vector(to_unsigned(scenario_full_18(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_18(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_18+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 19
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_19*2-1 loop
	assert RAM(SCENARIO_ADDRESS_19+i) = std_logic_vector(to_unsigned(scenario_full_19(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_19(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_19+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 20
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_20*2-1 loop
	assert RAM(SCENARIO_ADDRESS_20+i) = std_logic_vector(to_unsigned(scenario_full_20(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_20(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_20+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 21
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_21*2-1 loop
	assert RAM(SCENARIO_ADDRESS_21+i) = std_logic_vector(to_unsigned(scenario_full_21(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_21(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_21+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 22
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_22*2-1 loop
	assert RAM(SCENARIO_ADDRESS_22+i) = std_logic_vector(to_unsigned(scenario_full_22(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_22(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_22+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 23
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_23*2-1 loop
	assert RAM(SCENARIO_ADDRESS_23+i) = std_logic_vector(to_unsigned(scenario_full_23(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_23(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_23+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 24
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_24*2-1 loop
	assert RAM(SCENARIO_ADDRESS_24+i) = std_logic_vector(to_unsigned(scenario_full_24(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_24(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_24+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 25
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_25*2-1 loop
	assert RAM(SCENARIO_ADDRESS_25+i) = std_logic_vector(to_unsigned(scenario_full_25(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_25(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_25+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 26
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_26*2-1 loop
	assert RAM(SCENARIO_ADDRESS_26+i) = std_logic_vector(to_unsigned(scenario_full_26(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_26(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_26+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 27
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_27*2-1 loop
	assert RAM(SCENARIO_ADDRESS_27+i) = std_logic_vector(to_unsigned(scenario_full_27(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_27(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_27+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 28
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_28*2-1 loop
	assert RAM(SCENARIO_ADDRESS_28+i) = std_logic_vector(to_unsigned(scenario_full_28(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_28(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_28+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 29
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_29*2-1 loop
	assert RAM(SCENARIO_ADDRESS_29+i) = std_logic_vector(to_unsigned(scenario_full_29(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_29(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_29+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 30
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_30*2-1 loop
	assert RAM(SCENARIO_ADDRESS_30+i) = std_logic_vector(to_unsigned(scenario_full_30(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_30(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_30+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);


	--Scenario 31
	wait until rising_edge(tb_start);
	while tb_done /= '1' loop
		wait until rising_edge(tb_clk);
	end loop;

	assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

	for i in 0 to SCENARIO_LENGTH_31*2-1 loop
	assert RAM(SCENARIO_ADDRESS_31+i) = std_logic_vector(to_unsigned(scenario_full_31(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_31(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS_31+i)))) severity failure;
	end loop;

	wait until falling_edge(tb_start);
	assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
	wait until falling_edge(tb_done);

-- End Test

        assert false report "Simulation Ended! TEST PASSATO 8214" severity failure;
    end process;

end architecture;
